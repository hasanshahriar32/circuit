CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 39 227 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 41 167 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
961 0 0
2
5.90006e-315 5.26354e-315
0
13 Logic Switch~
5 574 244 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3178 0 0
2
5.90006e-315 5.30499e-315
0
13 Logic Switch~
5 575 147 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3409 0 0
2
5.90006e-315 5.32571e-315
0
13 Logic Switch~
5 289 156 0 1 11
0 17
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3951 0 0
2
5.90006e-315 5.34643e-315
0
13 Logic Switch~
5 288 253 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8885 0 0
2
5.90006e-315 5.3568e-315
0
14 Logic Display~
6 333 219 0 1 2
10 3
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
44498.5 0
0
14 Logic Display~
6 332 171 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
44498.5 0
0
7 Pulser~
4 117 403 0 10 12
0 7 2 5 2 0 0 15 15 8
7
0
0 0 4656 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 V
9442 0 0
2
44498.5 0
0
9 Inverter~
13 307 396 0 2 22
0 5 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9424 0 0
2
44498.5 1
0
2 +V
167 37 333 0 1 3
0 7
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9968 0 0
2
44498.5 2
0
7 Ground~
168 85 460 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9281 0 0
2
44498.5 3
0
14 Logic Display~
6 621 211 0 1 2
10 8
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
44498.5 4
0
14 Logic Display~
6 620 161 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
44498.5 5
0
14 Logic Display~
6 191 350 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
44498.5 6
0
9 2-In AND~
219 159 159 0 3 22
0 8 11 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4139 0 0
2
5.90006e-315 5.36716e-315
0
9 2-In AND~
219 160 238 0 3 22
0 10 9 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6435 0 0
2
5.90006e-315 5.37752e-315
0
5 4027~
219 575 215 0 7 32
0 15 4 6 3 14 8 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 1 0
1 U
5283 0 0
2
5.90006e-315 5.38788e-315
0
5 4027~
219 289 224 0 7 32
0 17 13 5 12 16 3 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
6874 0 0
2
44498.5 7
0
23
1 0 3 0 0 4096 0 7 0 0 18 2
333 205
333 206
1 0 4 0 0 4096 0 8 0 0 19 2
332 189
332 188
0 0 5 0 0 8192 0 0 0 7 5 4
190 394
190 391
231 391
231 396
2 3 6 0 0 4224 0 10 18 0 0 5
328 396
546 396
546 394
551 394
551 188
1 3 5 0 0 16512 0 10 19 0 0 6
292 396
231 396
231 394
233 394
233 197
265 197
1 1 7 0 0 8320 0 11 9 0 0 3
37 342
37 394
93 394
3 1 5 0 0 0 0 9 15 0 0 3
141 394
191 394
191 368
4 1 2 0 0 12416 0 9 12 0 0 5
147 403
151 403
151 441
85 441
85 454
2 1 2 0 0 0 0 9 12 0 0 5
87 403
83 403
83 446
85 446
85 454
1 0 8 0 0 0 0 13 0 0 14 2
621 197
621 197
1 0 9 0 0 0 0 14 0 0 15 2
620 179
620 179
1 1 10 0 0 4224 0 1 17 0 0 4
51 227
128 227
128 229
136 229
1 2 11 0 0 4224 0 2 16 0 0 4
53 167
127 167
127 168
135 168
6 1 8 0 0 12416 0 18 16 0 0 6
605 197
663 197
663 103
115 103
115 150
135 150
7 2 9 0 0 12416 0 18 17 0 0 6
599 179
639 179
639 284
117 284
117 247
136 247
3 4 12 0 0 4224 0 17 19 0 0 4
181 238
257 238
257 206
265 206
3 2 13 0 0 4224 0 16 19 0 0 4
180 159
257 159
257 188
265 188
6 4 3 0 0 4224 0 19 18 0 0 4
319 206
543 206
543 197
551 197
7 2 4 0 0 4224 0 19 18 0 0 4
313 188
543 188
543 179
551 179
1 5 14 0 0 4224 0 3 18 0 0 2
575 231
575 221
1 1 15 0 0 4224 0 4 18 0 0 2
575 159
575 158
1 5 16 0 0 4224 0 6 19 0 0 2
289 240
289 230
1 1 17 0 0 4224 0 5 19 0 0 2
289 168
289 167
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
53 149 76 173
60 154 68 170
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
50 213 73 237
57 218 65 234
1 K
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
39 67 182 91
46 73 174 89
16 Master Slave J-K
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
