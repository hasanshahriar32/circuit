CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 440 1364 717
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 417 88 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3171 0 0
2
44500.2 0
0
13 Logic Switch~
5 339 85 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4139 0 0
2
44500.2 0
0
13 Logic Switch~
5 268 90 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6435 0 0
2
44500.2 0
0
13 Logic Switch~
5 194 91 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
44500.2 0
0
6 74266~
219 487 421 0 3 22
0 13 3 11
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6874 0 0
2
44500.2 0
0
6 74266~
219 485 378 0 3 22
0 14 2 12
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5305 0 0
2
44500.2 0
0
14 Logic Display~
6 670 373 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
44500.2 0
0
14 Logic Display~
6 668 521 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
44500.2 0
0
14 Logic Display~
6 675 225 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
44500.2 0
0
9 2-In AND~
219 500 594 0 3 22
0 5 3 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3751 0 0
2
44500.2 0
0
8 3-In OR~
219 561 537 0 4 22
0 8 7 6 9
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
4292 0 0
2
44500.2 0
0
8 3-In OR~
219 559 242 0 4 22
0 18 17 16 15
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
6118 0 0
2
44500.2 0
0
9 2-In AND~
219 485 204 0 3 22
0 13 20 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
34 0 0
2
44500.2 0
0
5 7415~
219 497 548 0 4 22
0 4 3 2 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
6357 0 0
2
44500.2 0
0
5 7415~
219 496 498 0 4 22
0 5 4 2 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
319 0 0
2
44500.2 0
0
5 7415~
219 493 294 0 4 22
0 13 14 19 16
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
3976 0 0
2
44500.2 0
0
5 7415~
219 490 249 0 4 22
0 14 20 19 17
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
7634 0 0
2
44500.2 0
0
9 2-In AND~
219 577 394 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
523 0 0
2
44500.2 0
0
9 Inverter~
13 436 152 0 2 22
0 2 19
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6748 0 0
2
44500.2 0
0
9 Inverter~
13 379 151 0 2 22
0 3 20
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
6901 0 0
2
44500.2 0
0
9 Inverter~
13 301 157 0 2 22
0 14 4
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
842 0 0
2
44500.2 0
0
9 Inverter~
13 223 155 0 2 22
0 21 5
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3277 0 0
2
44500.2 0
0
43
3 0 2 0 0 4096 0 14 0 0 36 2
473 557
417 557
2 0 3 0 0 4096 0 14 0 0 38 2
473 548
339 548
1 0 4 0 0 4096 0 14 0 0 34 2
473 539
304 539
2 0 3 0 0 4096 0 10 0 0 38 2
476 603
339 603
1 0 5 0 0 4096 0 10 0 0 41 2
476 585
226 585
3 0 2 0 0 0 0 15 0 0 36 2
472 507
417 507
2 0 4 0 0 0 0 15 0 0 34 2
472 498
304 498
1 0 5 0 0 0 0 15 0 0 41 2
472 489
226 489
3 3 6 0 0 8320 0 11 10 0 0 4
548 546
535 546
535 594
521 594
2 4 7 0 0 4224 0 11 14 0 0 4
549 537
526 537
526 548
518 548
1 4 8 0 0 8320 0 11 15 0 0 4
548 528
524 528
524 498
517 498
4 1 9 0 0 8320 0 11 8 0 0 3
594 537
594 539
668 539
1 3 10 0 0 8320 0 7 18 0 0 3
670 391
670 394
598 394
2 3 11 0 0 8320 0 18 5 0 0 4
553 403
540 403
540 421
526 421
3 1 12 0 0 4224 0 6 18 0 0 4
524 378
540 378
540 385
553 385
2 0 3 0 0 0 0 5 0 0 38 2
471 430
339 430
1 0 13 0 0 4096 0 5 0 0 43 2
471 412
194 412
2 0 2 0 0 0 0 6 0 0 36 2
469 387
417 387
1 0 14 0 0 4096 0 6 0 0 40 2
469 369
268 369
1 4 15 0 0 8320 0 9 12 0 0 3
675 243
675 242
592 242
3 4 16 0 0 8320 0 12 16 0 0 4
546 251
532 251
532 294
514 294
2 4 17 0 0 4224 0 12 17 0 0 4
547 242
527 242
527 249
511 249
1 3 18 0 0 8320 0 12 13 0 0 4
546 233
525 233
525 204
506 204
3 0 19 0 0 4096 0 16 0 0 32 2
469 303
439 303
2 0 14 0 0 0 0 16 0 0 40 2
469 294
268 294
1 0 13 0 0 0 0 16 0 0 43 2
469 285
194 285
3 0 19 0 0 0 0 17 0 0 32 2
466 258
439 258
2 0 20 0 0 4096 0 17 0 0 33 2
466 249
382 249
1 0 14 0 0 0 0 17 0 0 40 2
466 240
268 240
2 0 20 0 0 0 0 13 0 0 33 2
461 213
382 213
1 0 13 0 0 0 0 13 0 0 43 2
461 195
194 195
2 0 19 0 0 4224 0 19 0 0 0 2
439 170
439 733
2 0 20 0 0 4224 0 20 0 0 0 2
382 169
382 733
2 0 4 0 0 4224 0 21 0 0 0 2
304 175
304 718
0 1 2 0 0 0 0 0 19 36 0 3
417 121
439 121
439 134
1 0 2 0 0 4224 0 1 0 0 0 3
417 100
417 702
420 702
0 1 3 0 0 0 0 0 20 38 0 3
339 122
382 122
382 133
1 0 3 0 0 4224 0 2 0 0 0 2
339 97
339 711
0 1 14 0 0 0 0 0 21 40 0 3
268 123
304 123
304 139
1 0 14 0 0 4224 0 3 0 0 0 3
268 102
268 673
271 673
2 0 5 0 0 4224 0 22 0 0 0 2
226 173
226 651
0 1 21 0 0 4224 0 0 22 0 0 3
197 118
226 118
226 137
1 0 13 0 0 4224 0 4 0 0 0 2
194 103
194 626
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
696 525 741 549
706 533 730 549
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
695 383 740 407
705 391 729 407
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
719 222 764 246
729 230 753 246
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
401 26 438 50
411 34 427 50
2 BO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
331 26 368 50
341 34 357 50
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
257 30 294 54
267 38 283 54
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
190 25 227 49
200 33 216 49
2 A1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
