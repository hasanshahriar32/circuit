CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 803 367 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44500.1 0
0
13 Logic Switch~
5 764 314 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44500.1 0
0
13 Logic Switch~
5 796 177 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44500.1 0
0
13 Logic Switch~
5 757 138 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
44500.1 0
0
13 Logic Switch~
5 123 502 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
44500.1 0
0
13 Logic Switch~
5 60 484 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
44500.1 0
0
13 Logic Switch~
5 117 372 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
44500.1 0
0
13 Logic Switch~
5 68 354 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
44500.1 0
0
13 Logic Switch~
5 86 214 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
44500.1 0
0
13 Logic Switch~
5 50 196 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
44500.1 0
0
13 Logic Switch~
5 82 133 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
44500.1 0
0
13 Logic Switch~
5 43 107 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9998 0 0
2
44500.1 0
0
14 Logic Display~
6 1250 189 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
44500.1 0
0
14 Logic Display~
6 558 389 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
44500.1 0
0
14 Logic Display~
6 432 130 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
44500.1 0
0
9 2-In NOR~
219 1142 222 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3670 0 0
2
44500.1 0
0
9 2-In NOR~
219 1026 329 0 3 22
0 5 3 6
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5616 0 0
2
44500.1 0
0
9 2-In NOR~
219 877 322 0 3 22
0 4 4 5
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
9323 0 0
2
44500.1 0
0
9 2-In NOR~
219 1027 164 0 3 22
0 9 8 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
317 0 0
2
44500.1 0
0
9 2-In NOR~
219 879 147 0 3 22
0 10 10 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3108 0 0
2
44500.1 0
0
10 2-In NAND~
219 435 427 0 3 22
0 16 15 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
44500.1 0
0
10 2-In NAND~
219 319 497 0 3 22
0 12 14 15
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
44500.1 0
0
10 2-In NAND~
219 207 515 0 3 22
0 13 13 14
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7876 0 0
2
44500.1 0
0
10 2-In NAND~
219 313 364 0 3 22
0 19 17 16
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6369 0 0
2
44500.1 0
0
10 2-In NAND~
219 203 378 0 3 22
0 18 18 17
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9172 0 0
2
44500.1 0
0
8 2-In OR~
219 324 157 0 3 22
0 21 22 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7100 0 0
2
44500.1 0
0
9 Inverter~
13 142 215 0 2 22
0 24 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3820 0 0
2
44500.1 0
0
9 2-In AND~
219 235 203 0 3 22
0 25 23 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7678 0 0
2
44500.1 0
0
9 Inverter~
13 141 129 0 2 22
0 27 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
961 0 0
2
44500.1 0
0
9 2-In AND~
219 228 118 0 3 22
0 28 26 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3178 0 0
2
44500.1 0
0
31
3 1 2 0 0 4224 0 16 13 0 0 3
1181 222
1250 222
1250 207
1 2 3 0 0 4224 0 1 17 0 0 4
815 367
1005 367
1005 338
1013 338
2 0 4 0 0 4096 0 18 0 0 4 3
864 331
834 331
834 314
1 1 4 0 0 4224 0 2 18 0 0 4
776 314
856 314
856 313
864 313
3 1 5 0 0 4224 0 18 17 0 0 4
916 322
1005 322
1005 320
1013 320
2 3 6 0 0 8320 0 16 17 0 0 4
1129 231
1073 231
1073 329
1065 329
3 1 7 0 0 4224 0 19 16 0 0 4
1066 164
1121 164
1121 213
1129 213
2 1 8 0 0 4224 0 19 3 0 0 4
1014 173
817 173
817 177
808 177
3 1 9 0 0 4224 0 20 19 0 0 4
918 147
1006 147
1006 155
1014 155
2 0 10 0 0 4096 0 20 0 0 11 3
866 156
841 156
841 138
1 1 10 0 0 4224 0 4 20 0 0 2
769 138
866 138
3 1 11 0 0 4224 0 21 14 0 0 3
462 427
558 427
558 407
1 1 12 0 0 4224 0 6 22 0 0 4
72 484
287 484
287 488
295 488
2 0 13 0 0 4096 0 23 0 0 15 3
183 524
148 524
148 502
1 1 13 0 0 4224 0 5 23 0 0 4
135 502
175 502
175 506
183 506
2 3 14 0 0 4224 0 22 23 0 0 4
295 506
242 506
242 515
234 515
3 2 15 0 0 8320 0 22 21 0 0 4
346 497
403 497
403 436
411 436
3 1 16 0 0 4224 0 24 21 0 0 4
340 364
403 364
403 418
411 418
3 2 17 0 0 4224 0 25 24 0 0 4
230 378
281 378
281 373
289 373
0 2 18 0 0 8192 0 0 25 21 0 3
148 372
148 387
179 387
1 1 18 0 0 4224 0 7 25 0 0 4
129 372
171 372
171 369
179 369
1 1 19 0 0 4224 0 8 24 0 0 4
80 354
281 354
281 355
289 355
3 1 20 0 0 4224 0 26 15 0 0 3
357 157
432 157
432 148
3 1 21 0 0 4224 0 30 26 0 0 4
249 118
303 118
303 148
311 148
3 2 22 0 0 4224 0 28 26 0 0 4
256 203
303 203
303 166
311 166
2 2 23 0 0 4224 0 27 28 0 0 4
163 215
203 215
203 212
211 212
1 1 24 0 0 4224 0 9 27 0 0 4
98 214
119 214
119 215
127 215
1 1 25 0 0 4224 0 10 28 0 0 4
62 196
203 196
203 194
211 194
2 2 26 0 0 4224 0 29 30 0 0 4
162 129
196 129
196 127
204 127
1 1 27 0 0 4224 0 11 29 0 0 4
94 133
118 133
118 129
126 129
1 1 28 0 0 4224 0 12 30 0 0 4
55 107
196 107
196 109
204 109
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
