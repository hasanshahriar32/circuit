CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 177 105 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44471.6 0
0
13 Logic Switch~
5 109 103 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44471.6 0
0
13 Logic Switch~
5 42 107 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44471.6 0
0
14 Logic Display~
6 872 117 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
44471.6 0
0
14 Logic Display~
6 954 114 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
44471.6 0
0
8 2-In OR~
219 722 353 0 3 22
0 7 6 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
44471.6 0
0
9 2-In AND~
219 608 238 0 3 22
0 3 8 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8901 0 0
2
44471.6 0
0
9 2-In AND~
219 333 263 0 3 22
0 2 9 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7361 0 0
2
44471.6 0
0
6 74136~
219 597 154 0 3 22
0 8 3 5
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
44471.6 0
0
6 74136~
219 325 178 0 3 22
0 9 2 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
44471.6 0
0
15
0 1 2 0 0 4096 0 0 8 11 0 3
276 187
276 254
309 254
0 1 3 0 0 4096 0 0 7 9 0 3
549 178
549 229
584 229
3 1 4 0 0 8320 0 6 4 0 0 3
755 353
872 353
872 135
3 1 5 0 0 4224 0 9 5 0 0 3
630 154
954 154
954 132
3 2 6 0 0 4224 0 8 6 0 0 4
354 263
696 263
696 362
709 362
3 1 7 0 0 8320 0 7 6 0 0 4
629 238
701 238
701 344
709 344
0 2 8 0 0 4096 0 0 7 8 0 3
515 145
515 247
584 247
0 1 8 0 0 4224 0 0 9 15 0 2
42 145
581 145
3 2 3 0 0 4224 0 10 9 0 0 4
358 178
568 178
568 163
581 163
0 2 9 0 0 4096 0 0 8 12 0 3
227 169
227 272
309 272
0 2 2 0 0 4096 0 0 10 13 0 2
177 187
309 187
0 1 9 0 0 4096 0 0 10 14 0 2
109 169
309 169
1 0 2 0 0 4224 0 1 0 0 0 2
177 117
177 436
1 0 9 0 0 4224 0 2 0 0 0 2
109 115
109 438
1 0 8 0 0 128 0 3 0 0 0 2
42 119
42 437
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
463 32 564 56
473 40 553 56
10 FULL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
841 68 902 92
851 76 891 92
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
931 65 976 89
941 73 965 89
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
98 40 123 64
106 48 114 64
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
162 42 191 66
172 50 180 66
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
29 39 58 63
39 47 47 63
1 X
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
