CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 50 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 365 121 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3978 0 0
2
5.90003e-315 0
0
13 Logic Switch~
5 208 125 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3494 0 0
2
5.90003e-315 5.26354e-315
0
13 Logic Switch~
5 50 129 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3507 0 0
2
5.90003e-315 0
0
5 7415~
219 651 530 0 4 22
0 5 6 3 11
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
5151 0 0
2
5.90003e-315 5.37752e-315
0
14 Logic Display~
6 786 522 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
5.90003e-315 5.36716e-315
0
14 Logic Display~
6 787 601 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8585 0 0
2
5.90003e-315 5.3568e-315
0
5 7415~
219 652 609 0 4 22
0 5 6 2 10
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
8809 0 0
2
5.90003e-315 5.34643e-315
0
5 7415~
219 651 773 0 4 22
0 5 4 2 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
5993 0 0
2
5.90003e-315 5.32571e-315
0
14 Logic Display~
6 786 765 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8654 0 0
2
5.90003e-315 5.30499e-315
0
14 Logic Display~
6 785 686 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7223 0 0
2
5.90003e-315 5.26354e-315
0
5 7415~
219 650 694 0 4 22
0 5 4 3 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
3641 0 0
2
5.90003e-315 0
0
5 7415~
219 650 380 0 4 22
0 7 4 3 13
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
3104 0 0
2
5.90003e-315 5.32571e-315
0
14 Logic Display~
6 785 372 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
5.90003e-315 5.30499e-315
0
14 Logic Display~
6 786 451 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
5.90003e-315 5.26354e-315
0
5 7415~
219 651 459 0 4 22
0 7 4 2 12
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
949 0 0
2
5.90003e-315 0
0
5 7415~
219 652 295 0 4 22
0 7 6 2 14
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
3371 0 0
2
5.90003e-315 5.26354e-315
0
14 Logic Display~
6 787 287 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7311 0 0
2
5.90003e-315 0
0
14 Logic Display~
6 786 208 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90003e-315 0
0
9 Inverter~
13 423 165 0 2 22
0 2 3
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
3526 0 0
2
5.90003e-315 5.26354e-315
0
9 Inverter~
13 266 169 0 2 22
0 4 6
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4129 0 0
2
5.90003e-315 0
0
9 Inverter~
13 108 175 0 2 22
0 5 7
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
6278 0 0
2
5.90003e-315 0
0
5 7415~
219 651 216 0 4 22
0 7 6 3 15
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3482 0 0
2
5.90003e-315 0
0
41
0 3 2 0 0 4096 0 0 8 35 0 2
365 782
627 782
0 3 3 0 0 4096 0 0 11 34 0 2
426 703
626 703
0 2 4 0 0 4096 0 0 8 38 0 2
208 773
627 773
0 2 4 0 0 0 0 0 11 38 0 2
208 694
626 694
0 1 5 0 0 4096 0 0 4 9 0 2
50 521
627 521
0 1 5 0 0 4096 0 0 7 9 0 2
50 600
628 600
0 1 5 0 0 0 0 0 11 9 0 2
50 685
626 685
0 1 5 0 0 0 0 0 8 9 0 2
50 764
627 764
0 0 5 0 0 4224 0 0 0 41 0 2
50 149
50 899
0 3 2 0 0 4096 0 0 7 35 0 2
365 618
628 618
0 2 6 0 0 4096 0 0 7 37 0 2
269 609
628 609
0 3 3 0 0 4096 0 0 4 34 0 2
426 539
627 539
0 2 6 0 0 0 0 0 4 37 0 2
269 530
627 530
0 3 2 0 0 0 0 0 15 35 0 2
365 468
627 468
0 2 4 0 0 0 0 0 15 38 0 2
208 459
627 459
0 1 7 0 0 4096 0 0 15 40 0 2
111 450
627 450
0 3 3 0 0 0 0 0 12 34 0 2
426 389
626 389
0 2 4 0 0 0 0 0 12 38 0 2
208 380
626 380
0 1 7 0 0 0 0 0 12 40 0 2
111 371
626 371
0 3 2 0 0 0 0 0 16 35 0 2
365 304
628 304
0 2 6 0 0 0 0 0 16 37 0 2
269 295
628 295
0 1 7 0 0 4096 0 0 16 40 0 2
111 286
628 286
0 3 3 0 0 0 0 0 22 34 0 2
426 225
627 225
0 2 6 0 0 0 0 0 22 37 0 2
269 216
627 216
0 1 7 0 0 0 0 0 22 40 0 2
111 207
627 207
4 1 8 0 0 4224 0 8 9 0 0 5
672 773
774 773
774 791
786 791
786 783
4 1 9 0 0 4224 0 11 10 0 0 5
671 694
773 694
773 712
785 712
785 704
4 1 10 0 0 4224 0 7 6 0 0 5
673 609
775 609
775 627
787 627
787 619
4 1 11 0 0 4224 0 4 5 0 0 5
672 530
774 530
774 548
786 548
786 540
4 1 12 0 0 4224 0 15 14 0 0 5
672 459
774 459
774 477
786 477
786 469
4 1 13 0 0 4224 0 12 13 0 0 5
671 380
773 380
773 398
785 398
785 390
4 1 14 0 0 4224 0 16 17 0 0 5
673 295
775 295
775 313
787 313
787 305
4 1 15 0 0 4224 0 22 18 0 0 5
672 216
774 216
774 234
786 234
786 226
2 0 3 0 0 4224 0 19 0 0 0 2
426 183
426 830
0 0 2 0 0 4224 0 0 0 36 0 2
365 141
365 896
1 1 2 0 0 0 0 1 19 0 0 4
365 133
365 141
426 141
426 147
2 0 6 0 0 4224 0 20 0 0 0 2
269 187
269 885
0 0 4 0 0 4224 0 0 0 39 0 2
208 145
208 894
1 1 4 0 0 0 0 2 20 0 0 4
208 137
208 145
269 145
269 151
2 0 7 0 0 4224 0 21 0 0 0 2
111 193
111 907
1 1 5 0 0 0 0 3 21 0 0 4
50 141
50 149
111 149
111 157
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
34 72 63 96
44 80 52 96
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
192 68 221 92
202 76 210 92
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
349 64 378 88
359 72 367 88
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 194 823 218
796 202 812 218
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
787 273 824 297
797 281 813 297
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 358 822 382
795 366 811 382
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 437 823 461
796 445 812 461
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 508 823 532
796 516 812 532
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
787 587 824 611
797 595 813 611
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 672 822 696
795 680 811 696
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 751 823 775
796 759 812 775
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
562 65 639 89
572 73 628 89
7 Decoder
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
