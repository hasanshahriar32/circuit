CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1534 620
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.240664 0.500000
176 629 1534 803
76546066 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 111 249 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
44500.3 0
0
9 2-In AND~
219 485 145 0 3 22
0 3 4 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9998 0 0
2
44500.3 0
0
5 SCOPE
12 354 403 0 1 11
0 7
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3536 0 0
2
44500.3 0
0
5 SCOPE
12 374 224 0 1 11
0 3
0
0 0 57584 0
2 Q1
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4597 0 0
2
44500.3 0
0
5 SCOPE
12 498 227 0 1 11
0 4
0
0 0 57584 0
2 Q2
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3835 0 0
2
44500.3 0
0
5 SCOPE
12 627 229 0 1 11
0 5
0
0 0 57584 0
2 Q3
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3670 0 0
2
44500.3 0
0
7 Ground~
168 192 501 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5616 0 0
2
44500.3 0
0
2 +V
167 107 400 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9323 0 0
2
44500.3 0
0
7 Pulser~
4 193 440 0 10 12
0 8 2 7 2 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
317 0 0
2
44500.3 0
0
14 Logic Display~
6 307 394 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
44500.3 0
0
14 Logic Display~
6 337 218 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
44500.3 0
0
14 Logic Display~
6 469 225 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
44500.3 0
0
14 Logic Display~
6 596 220 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
44500.3 0
0
5 4027~
219 537 310 0 7 32
0 11 6 7 6 12 13 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
6369 0 0
2
44500.3 0
0
5 4027~
219 412 307 0 7 32
0 14 3 7 3 15 16 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
9172 0 0
2
44500.3 0
0
5 4027~
219 267 307 0 7 32
0 17 10 7 10 18 19 3
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
7100 0 0
2
44500.3 0
0
25
1 0 3 0 0 4096 0 11 0 0 23 2
337 236
337 271
1 0 3 0 0 0 0 4 0 0 23 2
374 236
374 271
1 0 4 0 0 8192 0 5 0 0 22 4
498 239
498 266
448 266
448 271
1 0 4 0 0 0 0 12 0 0 22 3
469 243
469 247
448 247
1 0 5 0 0 8192 0 6 0 0 18 3
627 241
627 248
561 248
1 0 5 0 0 0 0 13 0 0 18 3
596 238
596 242
561 242
4 0 6 0 0 8192 0 14 0 0 20 3
513 292
508 292
508 264
0 4 3 0 0 0 0 0 15 23 0 3
364 271
364 289
388 289
0 3 7 0 0 4096 0 0 14 12 0 4
354 423
496 423
496 283
513 283
0 3 7 0 0 4224 0 0 15 12 0 3
342 426
342 280
388 280
1 0 7 0 0 0 0 10 0 0 12 2
307 412
307 426
1 0 7 0 0 0 0 3 0 0 13 3
354 415
354 426
254 426
3 3 7 0 0 0 0 9 16 0 0 6
217 431
254 431
254 384
185 384
185 280
243 280
1 0 2 0 0 4096 0 7 0 0 15 2
192 495
192 478
2 4 2 0 0 12416 0 9 9 0 0 6
163 440
152 440
152 478
242 478
242 440
223 440
1 1 8 0 0 8320 0 8 9 0 0 3
107 409
107 431
169 431
0 0 9 0 0 4224 0 0 0 0 0 2
640 149
649 149
7 0 5 0 0 4224 0 14 0 0 0 3
561 274
561 158
595 158
0 0 6 0 0 8192 0 0 0 20 0 3
518 145
518 140
595 140
3 2 6 0 0 8320 0 2 14 0 0 6
506 145
520 145
520 249
508 249
508 274
513 274
0 1 3 0 0 4224 0 0 2 23 0 3
382 271
382 136
461 136
7 2 4 0 0 8320 0 15 2 0 0 4
436 271
448 271
448 154
461 154
7 2 3 0 0 0 0 16 15 0 0 2
291 271
388 271
0 4 10 0 0 4096 0 0 16 25 0 3
207 249
207 289
243 289
1 2 10 0 0 4224 0 1 16 0 0 4
123 249
235 249
235 271
243 271
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
