CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 17 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
71 C:\Program Files (x86)\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
143654930 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 815 295 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44499.8 1
0
13 Logic Switch~
5 808 165 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44499.8 2
0
13 Logic Switch~
5 697 276 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44499.8 3
0
13 Logic Switch~
5 686 156 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44499.8 4
0
13 Logic Switch~
5 571 286 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44499.8 5
0
13 Logic Switch~
5 566 162 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44499.8 6
0
13 Logic Switch~
5 457 285 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44499.8 7
0
13 Logic Switch~
5 447 158 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44499.8 8
0
13 Logic Switch~
5 323 159 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44499.8 9
0
13 Logic Switch~
5 330 278 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
44499.8 10
0
13 Logic Switch~
5 229 98 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
44499.8 11
0
2 +V
167 178 275 0 1 3
0 9
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
44499.8 0
0
7 Ground~
168 215 396 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
44499.8 13
0
9 Inverter~
13 286 199 0 2 22
0 3 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 4 0
1 U
4597 0 0
2
44499.8 14
0
9 Inverter~
13 783 226 0 2 22
0 5 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 4 4 0
1 U
3835 0 0
2
44499.8 15
0
9 Inverter~
13 664 227 0 2 22
0 6 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 3 4 0
1 U
3670 0 0
2
44499.8 16
0
9 Inverter~
13 538 229 0 2 22
0 7 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 4 0
1 U
5616 0 0
2
44499.8 17
0
9 Inverter~
13 408 229 0 2 22
0 8 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 4 0
1 U
9323 0 0
2
44499.8 18
0
14 Logic Display~
6 992 396 0 1 2
10 27
0
0 0 53856 180
6 100MEG
3 -16 45 -8
3 L10
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44499.8 19
0
14 Logic Display~
6 761 399 0 1 2
10 20
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44499.8 20
0
14 Logic Display~
6 635 403 0 1 2
10 19
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44499.8 21
0
14 Logic Display~
6 508 403 0 1 2
10 28
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
44499.8 22
0
14 Logic Display~
6 387 404 0 1 2
10 22
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
44499.8 23
0
14 Logic Display~
6 751 67 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
44499.8 24
0
14 Logic Display~
6 625 67 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
44499.8 25
0
14 Logic Display~
6 510 67 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
44499.8 26
0
14 Logic Display~
6 395 67 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
44499.8 27
0
7 Pulser~
4 243 347 0 10 12
0 9 2 30 2 0 0 5 5 4
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 V
7678 0 0
2
44499.8 28
0
5 4027~
219 826 244 0 7 32
0 18 5 30 23 17 27 29
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 1 3 0
1 U
961 0 0
2
44499.8 29
0
5 4027~
219 707 245 0 7 32
0 15 6 30 24 16 20 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 2 2 0
1 U
3178 0 0
2
44499.8 30
0
5 4027~
219 582 247 0 7 32
0 14 7 30 25 13 19 6
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 1 2 0
1 U
3409 0 0
2
44499.8 31
0
5 4027~
219 465 245 0 7 32
0 12 8 30 21 11 28 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 2 1 0
1 U
3951 0 0
2
44499.8 32
0
5 4027~
219 350 242 0 7 32
0 10 3 30 4 26 22 8
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 1928712129
65 0 0 0 2 1 1 0
1 U
8885 0 0
2
44499.8 33
0
14 Logic Display~
6 988 178 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
44499.8 34
0
45
0 2 3 0 0 4096 0 0 33 10 0 4
263 185
317 185
317 206
326 206
2 4 4 0 0 8320 0 14 33 0 0 4
307 199
313 199
313 224
326 224
0 2 5 0 0 4096 0 0 29 36 0 2
751 209
802 208
0 2 6 0 0 4096 0 0 30 37 0 2
625 209
683 209
0 2 7 0 0 4096 0 0 31 38 0 4
509 183
550 183
550 211
558 211
0 2 8 0 0 4096 0 0 32 39 0 4
395 195
433 195
433 209
441 209
4 1 2 0 0 12416 0 28 13 0 0 5
273 347
277 347
277 382
215 382
215 390
2 1 2 0 0 0 0 28 13 0 0 5
213 347
209 347
209 382
215 382
215 390
1 1 9 0 0 20608 0 12 28 0 0 7
178 284
178 288
195 288
195 287
205 287
205 338
219 338
1 1 3 0 0 8320 0 11 14 0 0 4
241 98
263 98
263 199
271 199
1 1 10 0 0 4224 0 33 9 0 0 3
350 185
350 159
335 159
1 5 11 0 0 8320 0 7 32 0 0 5
469 285
474 285
474 259
465 259
465 251
1 1 12 0 0 4224 0 32 8 0 0 3
465 188
465 158
459 158
1 5 13 0 0 8320 0 5 31 0 0 5
583 286
588 286
588 261
582 261
582 253
1 1 14 0 0 8320 0 6 31 0 0 3
578 162
582 162
582 190
1 1 15 0 0 8320 0 4 30 0 0 3
698 156
707 156
707 188
5 1 16 0 0 4224 0 30 3 0 0 5
707 251
707 266
718 266
718 276
709 276
1 5 17 0 0 8320 0 1 29 0 0 5
827 295
832 295
832 258
826 258
826 250
1 1 18 0 0 8320 0 2 29 0 0 3
820 165
826 165
826 187
6 0 19 0 0 4096 0 31 0 0 33 2
612 229
634 229
6 1 20 0 0 8320 0 30 20 0 0 3
737 227
761 227
761 385
0 1 5 0 0 0 0 0 15 36 0 4
751 179
760 179
760 226
768 226
0 1 6 0 0 0 0 0 16 37 0 4
625 177
641 177
641 227
649 227
0 1 7 0 0 0 0 0 17 38 0 4
509 199
515 199
515 229
523 229
2 4 21 0 0 12416 0 18 32 0 0 4
429 229
433 229
433 227
441 227
6 1 22 0 0 8320 0 33 23 0 0 3
380 224
387 224
387 390
0 1 8 0 0 0 0 0 18 39 0 3
385 205
385 229
393 229
2 4 23 0 0 4224 0 15 29 0 0 2
804 226
802 226
2 4 24 0 0 4224 0 16 30 0 0 2
685 227
683 227
2 4 25 0 0 4224 0 17 31 0 0 2
559 229
558 229
5 1 26 0 0 4224 0 33 10 0 0 3
350 248
350 278
342 278
6 1 27 0 0 8320 0 29 19 0 0 3
856 226
992 226
992 382
0 1 19 0 0 4224 0 0 21 0 0 3
634 229
634 389
635 389
6 1 28 0 0 8320 0 32 22 0 0 3
495 227
508 227
508 389
7 1 29 0 0 4224 0 29 34 0 0 3
850 208
988 208
988 196
7 1 5 0 0 8320 0 30 24 0 0 3
731 209
751 209
751 85
7 1 6 0 0 8320 0 31 25 0 0 3
606 211
625 211
625 85
7 1 7 0 0 8320 0 32 26 0 0 4
489 209
509 209
509 85
510 85
7 1 8 0 0 12416 0 33 27 0 0 4
374 206
374 205
395 205
395 85
3 0 30 0 0 12288 0 29 0 0 41 4
802 217
741 217
741 311
616 311
3 0 30 0 0 0 0 30 0 0 42 4
683 218
616 218
616 311
499 311
3 0 30 0 0 0 0 31 0 0 44 5
558 220
499 220
499 311
431 311
431 316
0 3 30 0 0 0 0 0 31 44 0 5
433 316
433 256
550 256
550 220
558 220
0 3 30 0 0 4224 0 0 32 45 0 4
281 316
433 316
433 218
441 218
3 3 30 0 0 0 0 33 28 0 0 4
326 215
281 215
281 338
267 338
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
525020 1079360 100 100 0 0
0 0 0 0
63 66 224 136
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 0.01 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
