CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 660 30 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
24 E:\Circuit Maker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 413 61 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44501.5 0
0
13 Logic Switch~
5 297 65 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44501.5 0
0
13 Logic Switch~
5 200 66 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44501.5 0
0
13 Logic Switch~
5 106 74 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44501.5 0
0
14 Logic Display~
6 808 1026 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
44501.5 0
0
14 Logic Display~
6 812 497 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
44501.5 0
0
14 Logic Display~
6 809 975 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
44501.5 0
0
14 Logic Display~
6 812 910 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
44501.5 0
0
14 Logic Display~
6 818 854 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
44501.5 0
0
14 Logic Display~
6 818 789 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
44501.5 0
0
14 Logic Display~
6 819 731 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
44501.5 0
0
14 Logic Display~
6 816 662 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
44501.5 0
0
14 Logic Display~
6 815 591 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
44501.5 0
0
14 Logic Display~
6 807 540 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
44501.5 0
0
14 Logic Display~
6 812 432 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
44501.5 0
0
14 Logic Display~
6 812 377 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
44501.5 0
0
14 Logic Display~
6 809 308 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
44501.5 0
0
14 Logic Display~
6 808 254 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
44501.5 0
0
14 Logic Display~
6 809 188 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
317 0 0
2
44501.5 0
0
14 Logic Display~
6 807 123 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3108 0 0
2
44501.5 0
0
9 Inverter~
13 454 116 0 2 22
0 3 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
4299 0 0
2
44501.5 0
0
9 Inverter~
13 343 120 0 2 22
0 24 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
9672 0 0
2
44501.5 0
0
9 Inverter~
13 238 121 0 2 22
0 25 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
7876 0 0
2
44501.5 0
0
9 Inverter~
13 148 135 0 2 22
0 8 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 9 0
1 U
6369 0 0
2
44501.5 0
0
9 4-In AND~
219 621 1038 0 5 22
0 8 25 24 3 7
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 8 0
1 U
9172 0 0
2
44501.5 0
0
9 4-In AND~
219 608 982 0 5 22
0 8 25 24 5 13
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U8A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 8 0
1 U
7100 0 0
2
44501.5 0
0
9 4-In AND~
219 607 921 0 5 22
0 8 25 4 3 14
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U7B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
3820 0 0
2
44501.5 0
0
9 4-In AND~
219 610 867 0 5 22
0 8 25 4 5 15
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U7A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
7678 0 0
2
44501.5 0
0
9 4-In AND~
219 603 746 0 5 22
0 8 11 24 5 17
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U6B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 6 0
1 U
961 0 0
2
44501.5 0
0
9 4-In AND~
219 604 683 0 5 22
0 8 11 4 3 18
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U6A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 6 0
1 U
3178 0 0
2
44501.5 0
0
9 4-In AND~
219 607 807 0 5 22
0 8 11 24 3 16
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U5B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
3409 0 0
2
44501.5 0
0
9 4-In AND~
219 606 619 0 5 22
0 8 11 4 5 12
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U5A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3951 0 0
2
44501.5 0
0
9 4-In AND~
219 609 559 0 5 22
0 2 25 24 3 6
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 4 0
1 U
8885 0 0
2
44501.5 0
0
9 4-In AND~
219 609 503 0 5 22
0 2 25 24 5 9
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U4A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
3780 0 0
2
44501.5 0
0
9 4-In AND~
219 597 443 0 5 22
0 2 25 4 3 19
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 3 0
1 U
9265 0 0
2
44501.5 0
0
9 4-In AND~
219 599 398 0 5 22
0 2 25 4 5 10
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
9442 0 0
2
44501.5 0
0
9 4-In AND~
219 592 334 0 5 22
0 2 11 24 3 20
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
9424 0 0
2
44501.5 0
0
9 4-In AND~
219 591 270 0 5 22
0 2 11 24 5 22
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
9968 0 0
2
44501.5 0
0
9 4-In AND~
219 591 200 0 5 22
0 2 11 4 3 21
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
9281 0 0
2
44501.5 0
0
9 4-In AND~
219 590 146 0 5 22
0 2 11 4 5 23
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 1 0
1 U
8464 0 0
2
44501.5 0
0
94
1 0 2 0 0 4096 0 40 0 0 92 4
566 133
183 133
183 149
169 149
4 0 3 0 0 4096 0 27 0 0 85 2
583 935
413 935
3 0 4 0 0 4096 0 27 0 0 86 2
583 926
364 926
4 0 5 0 0 4096 0 26 0 0 83 2
584 996
475 996
5 1 6 0 0 8320 0 33 14 0 0 3
630 559
630 558
807 558
4 0 5 0 0 0 0 34 0 0 56 2
585 517
585 517
5 1 7 0 0 4224 0 25 5 0 0 5
642 1038
778 1038
778 1060
808 1060
808 1044
1 0 8 0 0 4096 0 25 0 0 94 2
597 1025
106 1025
5 1 9 0 0 4224 0 34 6 0 0 4
630 503
755 503
755 515
812 515
5 1 10 0 0 4224 0 36 16 0 0 3
620 398
812 398
812 395
2 0 11 0 0 4096 0 31 0 0 89 2
583 803
259 803
1 0 8 0 0 0 0 28 0 0 94 2
586 854
106 854
1 5 12 0 0 8320 0 13 32 0 0 3
815 609
815 619
627 619
5 1 13 0 0 4224 0 26 7 0 0 5
629 982
769 982
769 996
809 996
809 993
5 1 14 0 0 4224 0 27 8 0 0 5
628 921
755 921
755 937
812 937
812 928
5 1 15 0 0 8320 0 28 9 0 0 3
631 867
631 872
818 872
5 1 16 0 0 4224 0 31 10 0 0 2
628 807
818 807
5 1 17 0 0 8320 0 29 11 0 0 3
624 746
624 749
819 749
5 1 18 0 0 4224 0 30 12 0 0 3
625 683
816 683
816 680
5 1 19 0 0 4224 0 35 15 0 0 4
618 443
754 443
754 450
812 450
5 1 20 0 0 4224 0 37 17 0 0 3
613 334
809 334
809 326
5 1 21 0 0 4224 0 39 19 0 0 5
612 200
734 200
734 209
809 209
809 206
1 0 22 0 0 4096 0 18 0 0 0 2
808 272
808 263
5 1 22 0 0 8320 0 38 18 0 0 3
612 270
612 272
808 272
1 5 23 0 0 8320 0 20 40 0 0 3
807 141
807 146
611 146
4 0 3 0 0 4096 0 25 0 0 85 2
597 1052
413 1052
3 0 24 0 0 4096 0 25 0 0 88 2
597 1043
297 1043
2 0 25 0 0 4096 0 25 0 0 91 2
597 1034
200 1034
3 0 24 0 0 0 0 26 0 0 88 2
584 987
297 987
2 0 25 0 0 0 0 26 0 0 91 2
584 978
200 978
1 0 8 0 0 0 0 26 0 0 94 2
584 969
106 969
2 0 25 0 0 0 0 27 0 0 91 2
583 917
200 917
1 0 8 0 0 0 0 27 0 0 94 2
583 908
106 908
4 0 5 0 0 4096 0 28 0 0 83 2
586 881
475 881
3 0 4 0 0 4096 0 28 0 0 86 2
586 872
364 872
2 0 25 0 0 0 0 28 0 0 91 2
586 863
200 863
4 0 3 0 0 0 0 31 0 0 85 2
583 821
413 821
3 0 24 0 0 0 0 31 0 0 88 2
583 812
297 812
1 0 8 0 0 0 0 31 0 0 94 2
583 794
106 794
4 0 5 0 0 0 0 29 0 0 83 2
579 760
475 760
3 0 24 0 0 0 0 29 0 0 88 2
579 751
297 751
2 0 11 0 0 0 0 29 0 0 89 2
579 742
259 742
1 0 8 0 0 0 0 29 0 0 94 2
579 733
106 733
4 0 3 0 0 0 0 30 0 0 85 2
580 697
413 697
3 0 4 0 0 0 0 30 0 0 86 2
580 688
364 688
2 0 11 0 0 0 0 30 0 0 89 2
580 679
259 679
1 0 8 0 0 0 0 30 0 0 94 2
580 670
106 670
4 0 5 0 0 0 0 32 0 0 83 2
582 633
475 633
3 0 4 0 0 0 0 32 0 0 86 2
582 624
364 624
2 0 11 0 0 0 0 32 0 0 89 2
582 615
259 615
1 0 8 0 0 0 0 32 0 0 94 2
582 606
106 606
4 0 3 0 0 0 0 33 0 0 85 2
585 573
413 573
3 0 24 0 0 0 0 33 0 0 88 2
585 564
297 564
2 0 25 0 0 0 0 33 0 0 91 2
585 555
200 555
1 0 2 0 0 4096 0 33 0 0 92 2
585 546
169 546
0 0 5 0 0 4096 0 0 0 0 83 2
589 517
475 517
3 0 24 0 0 0 0 34 0 0 88 2
585 508
297 508
2 0 25 0 0 0 0 34 0 0 91 2
585 499
200 499
1 0 2 0 0 0 0 34 0 0 92 2
585 490
169 490
4 0 3 0 0 0 0 35 0 0 85 2
573 457
413 457
3 0 4 0 0 0 0 35 0 0 86 2
573 448
364 448
2 0 25 0 0 0 0 35 0 0 91 2
573 439
200 439
1 0 2 0 0 0 0 35 0 0 92 2
573 430
169 430
4 0 5 0 0 0 0 36 0 0 83 2
575 412
475 412
3 0 4 0 0 0 0 36 0 0 86 2
575 403
364 403
2 0 25 0 0 0 0 36 0 0 91 2
575 394
200 394
1 0 2 0 0 0 0 36 0 0 92 2
575 385
169 385
4 0 3 0 0 0 0 37 0 0 85 2
568 348
413 348
3 0 24 0 0 0 0 37 0 0 88 2
568 339
297 339
2 0 11 0 0 0 0 37 0 0 89 2
568 330
259 330
1 0 2 0 0 0 0 37 0 0 92 2
568 321
169 321
4 0 5 0 0 0 0 38 0 0 83 2
567 284
475 284
3 0 24 0 0 0 0 38 0 0 88 2
567 275
297 275
2 0 11 0 0 0 0 38 0 0 89 2
567 266
259 266
1 0 2 0 0 0 0 38 0 0 92 2
567 257
169 257
4 0 3 0 0 0 0 39 0 0 85 2
567 214
413 214
3 0 4 0 0 0 0 39 0 0 86 2
567 205
364 205
2 0 11 0 0 0 0 39 0 0 89 2
567 196
259 196
1 0 2 0 0 0 0 39 0 0 92 2
567 187
169 187
4 0 5 0 0 0 0 40 0 0 83 2
566 160
475 160
3 0 4 0 0 0 0 40 0 0 86 2
566 151
364 151
2 0 11 0 0 0 0 40 0 0 89 2
566 142
259 142
2 0 5 0 0 4224 0 21 0 0 0 2
475 116
475 1087
1 0 3 0 0 0 0 21 0 0 85 2
439 116
413 116
1 0 3 0 0 4224 0 1 0 0 0 2
413 73
413 1086
2 0 4 0 0 4224 0 22 0 0 0 2
364 120
364 1089
1 0 24 0 0 0 0 22 0 0 88 2
328 120
297 120
1 0 24 0 0 4224 0 2 0 0 0 2
297 77
297 1090
2 0 11 0 0 4224 0 23 0 0 0 2
259 121
259 1091
1 0 25 0 0 0 0 23 0 0 91 2
223 121
200 121
1 0 25 0 0 4224 0 3 0 0 0 2
200 78
200 1089
2 0 2 0 0 4224 0 24 0 0 0 2
169 135
169 1091
1 0 8 0 0 0 0 24 0 0 94 2
133 135
106 135
1 0 8 0 0 4224 0 4 0 0 0 2
106 86
106 1089
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
286 6 315 30
296 14 304 30
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
198 7 227 31
208 15 216 31
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
407 3 436 27
417 11 425 27
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
96 10 125 34
106 18 114 34
1 E
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
