CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9961490 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 527 148 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 1V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44656 4
0
13 Logic Switch~
5 359 366 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
3 -1V
-9 -16 12 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
44656 3
0
13 Logic Switch~
5 355 317 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
3 -1V
-9 -16 12 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
44656 2
0
13 Logic Switch~
5 356 266 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
3421 0 0
2
44656 1
0
13 Logic Switch~
5 353 220 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
8157 0 0
2
44656 0
0
7 Op Amp~
219 596 293 0 3 7
0 2 4 3
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
5572 0 0
2
44656 8
0
7 Ground~
168 559 338 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8901 0 0
2
44656 7
0
11 Multimeter~
205 773 257 0 21 21
0 3 10 11 2 0 0 0 0 0
32 51 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
1 R
7361 0 0
2
44656 6
0
7 Ground~
168 798 316 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4747 0 0
2
44656 5
0
9 Resistor~
219 625 230 0 2 5
0 4 3
0
0 0 880 0
1 8
-4 -14 3 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
972 0 0
2
44656 14
0
9 Resistor~
219 527 205 0 2 5
0 12 5
0
0 0 880 90
1 1
11 0 18 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 0 0 0 0
1 R
3472 0 0
2
44656 13
0
9 Resistor~
219 426 366 0 2 5
0 6 4
0
0 0 880 0
1 8
-4 -14 3 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9998 0 0
2
44656 12
0
9 Resistor~
219 421 317 0 2 5
0 7 4
0
0 0 880 0
1 4
-4 -14 3 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3536 0 0
2
44656 11
0
9 Resistor~
219 421 266 0 2 5
0 8 4
0
0 0 880 0
1 2
-4 -14 3 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4597 0 0
2
44656 10
0
9 Resistor~
219 423 220 0 2 5
0 9 4
0
0 0 880 0
1 1
-4 -14 3 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3835 0 0
2
44656 9
0
15
1 0 0 0 0 0 0 11 0 0 8 2
527 223
527 287
2 0 3 0 0 8208 0 10 0 0 4 3
643 230
673 230
673 293
1 4 2 0 0 4112 0 9 8 0 0 2
798 310
798 280
3 1 3 0 0 4240 0 6 8 0 0 3
614 293
748 293
748 280
1 0 4 0 0 8208 0 10 0 0 8 3
607 230
559 230
559 287
1 1 2 0 0 4240 0 7 6 0 0 3
559 332
559 299
578 299
1 2 5 0 0 4240 0 1 11 0 0 2
527 160
527 187
2 0 4 0 0 4112 0 6 0 0 15 2
578 287
479 287
1 1 6 0 0 4240 0 2 12 0 0 2
371 366
408 366
1 1 7 0 0 4240 0 3 13 0 0 2
367 317
403 317
1 1 8 0 0 4240 0 4 14 0 0 4
368 266
404 266
404 266
403 266
1 1 9 0 0 4240 0 5 15 0 0 4
365 220
406 220
406 220
405 220
2 0 4 0 0 16 0 13 0 0 15 2
439 317
479 317
2 0 4 0 0 16 0 14 0 0 15 2
439 266
479 266
2 2 4 0 0 8336 0 15 12 0 0 4
441 220
479 220
479 366
444 366
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
