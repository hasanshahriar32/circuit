CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 502
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.312600 0.500000
176 511 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 212 116 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
5.90027e-315 0
0
13 Logic Switch~
5 221 290 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6263 0 0
2
5.90027e-315 0
0
13 Logic Switch~
5 218 166 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
5.90027e-315 0
0
5 SCOPE
12 294 135 0 1 11
0 3
0
0 0 57584 270
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8783 0 0
2
44664.5 0
0
5 SCOPE
12 431 134 0 1 11
0 4
0
0 0 57584 270
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3221 0 0
2
44664.5 0
0
5 SCOPE
12 549 135 0 1 11
0 5
0
0 0 57584 270
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3215 0 0
2
44664.5 0
0
5 SCOPE
12 667 135 0 1 11
0 6
0
0 0 57584 270
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7903 0 0
2
44664.5 0
0
5 SCOPE
12 783 145 0 1 11
0 7
0
0 0 57584 270
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7121 0 0
2
44664.5 0
0
7 Pulser~
4 828 221 0 10 12
0 8 2 7 2 0 0 5 5 2
7
0
0 0 4656 180
0
2 V4
-7 -29 7 -21
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
4484 0 0
2
44664.4 0
0
2 +V
167 899 157 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5996 0 0
2
5.90027e-315 0
0
7 Ground~
168 825 265 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7804 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 287 77 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 422 78 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 540 77 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 659 82 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 775 80 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.90027e-315 0
0
6 74112~
219 337 255 0 7 32
0 10 9 4 9 11 12 3
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U2B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
7849 0 0
2
5.90027e-315 0
0
6 74112~
219 464 255 0 7 32
0 10 9 5 9 11 13 4
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U2A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
6343 0 0
2
5.90027e-315 0
0
6 74112~
219 584 255 0 7 32
0 10 9 6 9 11 14 5
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U1B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7376 0 0
2
5.90027e-315 0
0
6 74112~
219 702 255 0 7 32
0 10 9 7 9 11 15 6
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U1A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
9156 0 0
2
5.90027e-315 0
0
33
1 0 3 0 0 4096 0 4 0 0 14 2
285 138
287 138
1 0 4 0 0 0 0 5 0 0 13 2
422 137
422 137
1 0 5 0 0 0 0 6 0 0 12 2
540 138
540 138
1 0 6 0 0 4096 0 7 0 0 11 2
658 138
659 138
1 0 7 0 0 4096 0 8 0 0 6 2
774 148
775 148
0 1 7 0 0 4224 0 0 16 10 0 2
775 228
775 98
1 0 2 0 0 0 0 11 0 0 8 2
825 259
825 259
4 2 2 0 0 12416 0 9 9 0 0 6
798 219
786 219
786 259
867 259
867 219
858 219
1 1 8 0 0 8320 0 9 10 0 0 3
852 228
899 228
899 166
3 3 7 0 0 0 0 20 9 0 0 2
732 228
804 228
1 0 6 0 0 4224 0 15 0 0 31 2
659 100
659 237
1 0 5 0 0 4224 0 14 0 0 32 2
540 95
540 237
1 0 4 0 0 4224 0 13 0 0 33 2
422 96
422 237
1 7 3 0 0 4224 0 12 17 0 0 3
287 95
287 237
313 237
4 0 9 0 0 4096 0 17 0 0 16 2
361 219
388 219
2 0 9 0 0 8192 0 17 0 0 22 3
361 237
388 237
388 116
4 0 9 0 0 0 0 18 0 0 18 2
488 219
512 219
2 0 9 0 0 0 0 18 0 0 22 3
488 237
512 237
512 116
4 0 9 0 0 0 0 19 0 0 20 2
608 219
629 219
2 0 9 0 0 0 0 19 0 0 22 3
608 237
629 237
629 116
4 0 9 0 0 0 0 20 0 0 22 2
726 219
762 219
1 2 9 0 0 4224 0 1 20 0 0 4
224 116
762 116
762 237
726 237
1 0 10 0 0 4096 0 17 0 0 26 2
337 264
337 290
1 0 10 0 0 0 0 18 0 0 26 2
464 264
464 290
1 0 10 0 0 0 0 19 0 0 26 2
584 264
584 290
1 1 10 0 0 4224 0 2 20 0 0 3
233 290
702 290
702 264
5 0 11 0 0 4096 0 17 0 0 30 2
337 189
337 166
5 0 11 0 0 0 0 18 0 0 30 2
464 189
464 166
5 0 11 0 0 0 0 19 0 0 30 2
584 189
584 166
1 5 11 0 0 4224 0 3 20 0 0 3
230 166
702 166
702 189
3 7 6 0 0 0 0 19 20 0 0 4
614 228
646 228
646 237
678 237
3 7 5 0 0 0 0 18 19 0 0 4
494 228
529 228
529 237
560 237
3 7 4 0 0 0 0 17 18 0 0 4
367 228
402 228
402 237
440 237
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
