CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 1 100 10
176 80 1364 472
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.360447 0.500000
176 481 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 622 290 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
44664.4 0
0
13 Logic Switch~
5 245 135 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
44664.4 0
0
5 SCOPE
12 628 210 0 1 11
0 4
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3124 0 0
2
44664.4 0
0
5 SCOPE
12 513 216 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3421 0 0
2
44664.4 0
0
5 SCOPE
12 394 221 0 1 11
0 6
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8157 0 0
2
44664.4 0
0
5 SCOPE
12 267 231 0 1 11
0 7
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5572 0 0
2
44664.4 0
0
14 Logic Display~
6 385 178 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
44664.4 0
0
14 Logic Display~
6 253 180 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
44664.4 0
0
14 Logic Display~
6 502 180 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
44664.4 0
0
14 Logic Display~
6 658 177 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
44664.4 0
0
2 +V
167 127 209 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3472 0 0
2
44664.4 0
0
7 Ground~
168 212 302 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9998 0 0
2
44664.4 0
0
7 Pulser~
4 213 250 0 10 12
0 8 2 7 2 0 0 5 5 4
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
3536 0 0
2
44664.4 0
0
6 JK RN~
219 584 237 0 6 22
0 9 5 9 3 10 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
4597 0 0
2
44664.4 0
0
6 JK RN~
219 469 244 0 6 22
0 9 6 9 3 11 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
3835 0 0
2
44664.4 0
0
6 JK RN~
219 343 249 0 6 22
0 9 7 9 3 12 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
3670 0 0
2
44664.4 0
0
24
1 0 3 0 0 4096 0 1 0 0 8 2
622 302
622 301
1 0 4 0 0 4096 0 3 0 0 9 2
628 222
628 220
1 0 5 0 0 4096 0 4 0 0 17 2
513 228
513 227
1 0 6 0 0 4096 0 5 0 0 18 2
394 233
394 232
1 0 7 0 0 4096 0 6 0 0 16 2
267 243
267 241
4 0 3 0 0 4096 0 15 0 0 8 2
469 275
469 301
4 0 3 0 0 4096 0 14 0 0 8 2
584 268
584 301
4 0 3 0 0 8320 0 16 0 0 0 3
343 280
343 301
651 301
1 6 4 0 0 8320 0 10 14 0 0 3
658 195
658 220
608 220
1 0 5 0 0 4224 0 9 0 0 17 2
502 198
502 227
1 0 6 0 0 4224 0 7 0 0 18 2
385 196
385 232
1 0 7 0 0 4096 0 8 0 0 16 2
253 198
253 241
1 1 8 0 0 8320 0 11 13 0 0 3
127 218
127 241
189 241
1 0 2 0 0 0 0 12 0 0 15 2
212 296
212 296
4 2 2 0 0 8320 0 13 13 0 0 4
243 250
243 296
183 296
183 250
3 2 7 0 0 4224 0 13 16 0 0 2
237 241
312 241
6 2 5 0 0 0 0 15 14 0 0 6
493 227
519 227
519 255
547 255
547 229
553 229
6 2 6 0 0 0 0 16 15 0 0 6
367 232
402 232
402 265
429 265
429 236
438 236
1 0 9 0 0 4096 0 16 0 0 20 2
319 232
292 232
3 0 9 0 0 8192 0 16 0 0 24 3
319 250
292 250
292 135
1 0 9 0 0 0 0 15 0 0 22 2
445 227
420 227
3 0 9 0 0 0 0 15 0 0 24 3
445 245
420 245
420 135
1 0 9 0 0 0 0 14 0 0 24 2
560 220
544 220
1 3 9 0 0 4224 0 2 14 0 0 4
257 135
544 135
544 238
560 238
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
