CircuitMaker Text
5.6
Probes: 2
Q1_3
Transient Analysis
0 283 139 65280
U1_6
Operating Point
0 577 138 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 817 553
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.317125 0.500000
344 176 985 326
9961490 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 318 235 0 1 11
0 5
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8748 0 0
2
44661.6 0
0
13 Logic Switch~
5 243 236 0 1 11
0 6
0
0 0 21360 90
2 0V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7168 0 0
2
44661.6 0
0
13 Logic Switch~
5 174 239 0 1 11
0 7
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
631 0 0
2
44661.6 0
0
13 Logic Switch~
5 102 238 0 1 11
0 8
0
0 0 21360 90
2 0V
16 0 30 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9466 0 0
2
44661.6 0
0
2 +V
167 400 24 0 1 3
0 4
0
0 0 54256 0
1 8
-4 -22 3 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3266 0 0
2
44661.6 0
0
7 Ground~
168 55 218 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7693 0 0
2
44661.6 0
0
7 Op Amp~
219 459 137 0 3 7
0 2 3 13
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
3723 0 0
2
44661.6 0
0
7 Ground~
168 424 176 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3440 0 0
2
44661.6 0
0
9 Resistor~
219 401 77 0 3 5
0 4 3 1
0
0 0 880 270
1 3
14 0 21 8
3 R11
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6263 0 0
2
44661.6 0
0
9 Resistor~
219 54 175 0 3 5
0 2 9 -1
0
0 0 880 90
1 2
11 0 18 8
3 R10
7 -12 28 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4900 0 0
2
44661.6 0
0
9 Resistor~
219 138 132 0 2 5
0 10 9
0
0 0 880 180
1 1
-4 -14 3 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8783 0 0
2
44661.6 0
0
9 Resistor~
219 212 133 0 2 5
0 11 10
0
0 0 880 180
1 1
-4 -14 3 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3221 0 0
2
44661.6 0
0
9 Resistor~
219 282 132 0 2 5
0 12 11
0
0 0 880 180
1 1
-4 -14 3 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3215 0 0
2
44661.6 0
0
9 Resistor~
219 514 91 0 2 5
0 13 3
0
0 0 880 180
1 3
-4 -14 3 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7903 0 0
2
44661.6 0
0
9 Resistor~
219 104 175 0 2 5
0 8 9
0
0 0 880 90
1 2
11 0 18 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7121 0 0
2
44661.6 0
0
9 Resistor~
219 175 176 0 2 5
0 7 10
0
0 0 880 90
1 2
11 0 18 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4484 0 0
2
44661.6 0
0
9 Resistor~
219 244 181 0 2 5
0 6 11
0
0 0 880 90
1 2
11 0 18 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5996 0 0
2
44661.6 0
0
9 Resistor~
219 321 180 0 2 5
0 5 12
0
0 0 880 90
1 2
11 0 18 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7804 0 0
2
44661.6 0
0
9 Resistor~
219 378 132 0 2 5
0 12 3
0
0 0 880 0
1 2
-4 -14 3 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5523 0 0
2
44661.6 0
0
20
2 0 3 0 0 4096 0 9 0 0 20 2
401 95
401 131
1 1 4 0 0 8320 0 5 9 0 0 3
400 33
401 33
401 59
1 1 5 0 0 8320 0 1 18 0 0 3
319 222
321 222
321 198
1 1 6 0 0 4224 0 2 17 0 0 2
244 223
244 199
1 1 7 0 0 4224 0 3 16 0 0 2
175 226
175 194
1 1 8 0 0 8320 0 4 15 0 0 3
103 225
104 225
104 193
1 1 2 0 0 8192 0 10 6 0 0 3
54 193
55 193
55 212
2 0 9 0 0 4096 0 15 0 0 15 2
104 157
104 132
2 0 10 0 0 4096 0 16 0 0 14 2
175 158
175 133
2 0 11 0 0 4096 0 17 0 0 13 2
244 163
244 132
2 0 12 0 0 4096 0 18 0 0 12 2
321 162
321 132
1 1 12 0 0 4224 0 13 19 0 0 2
300 132
360 132
1 2 11 0 0 8320 0 12 13 0 0 3
230 133
230 132
264 132
1 2 10 0 0 8320 0 11 12 0 0 3
156 132
156 133
194 133
2 2 9 0 0 8320 0 10 11 0 0 3
54 157
54 132
120 132
1 1 2 0 0 8320 0 7 8 0 0 3
441 143
424 143
424 170
1 0 13 0 0 8192 0 14 0 0 18 3
532 91
555 91
555 137
3 0 13 0 0 4224 0 7 0 0 0 2
477 137
598 137
0 2 3 0 0 8320 0 0 14 20 0 3
416 131
416 91
496 91
2 2 3 0 0 0 0 19 7 0 0 3
396 132
396 131
441 131
0
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
