CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 210 1 110 10
165 80 1534 485
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
10 D:\BOM.DAT
0 7
5 2 0.435198 0.500000
165 494 1534 813
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 430 333 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 180
2 5V
-7 -16 7 -8
2 V3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3171 0 0
2
44499.6 0
0
5 SCOPE
12 112 391 0 1 11
0 3
0
0 0 57584 0
3 TP5
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4139 0 0
2
44499.6 0
0
5 SCOPE
12 153 410 0 1 11
0 4
0
0 0 57584 90
3 TP4
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6435 0 0
2
44499.6 0
0
5 SCOPE
12 227 409 0 1 11
0 5
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5283 0 0
2
44499.6 0
0
5 SCOPE
12 297 419 0 1 11
0 6
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6874 0 0
2
44499.6 0
0
5 SCOPE
12 399 385 0 1 11
0 7
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5305 0 0
2
44499.6 0
0
2 +V
167 355 487 0 1 3
0 9
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
34 0 0
2
44499.6 0
0
7 Ground~
168 394 542 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
969 0 0
2
44499.6 0
0
14 Logic Display~
6 236 446 0 1 2
10 6
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
44499.6 0
0
14 Logic Display~
6 199 446 0 1 2
10 5
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
44499.6 0
0
14 Logic Display~
6 164 445 0 1 2
10 4
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
44499.6 0
0
14 Logic Display~
6 126 445 0 1 2
10 3
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
44499.6 0
0
5 4081~
219 196 246 0 3 22
0 11 4 10
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
34 0 0
2
44499.6 0
0
5 4081~
219 272 249 0 3 22
0 6 5 11
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6357 0 0
2
44499.6 0
0
7 Pulser~
4 385 507 0 10 12
0 9 2 7 2 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
319 0 0
2
44499.6 0
0
5 4027~
219 340 361 0 7 32
0 12 8 7 8 13 14 6
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3976 0 0
2
44499.6 0
0
5 4027~
219 117 358 0 7 32
0 15 10 7 10 16 17 3
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U2A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7634 0 0
2
44499.6 0
0
5 4027~
219 193 359 0 7 32
0 18 11 7 11 19 20 4
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U1B
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
523 0 0
2
44499.6 0
0
5 4027~
219 270 361 0 7 32
0 21 6 7 6 22 23 5
0
0 0 4720 512
4 4027
7 -60 35 -52
3 U1A
27 -61 48 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6748 0 0
2
44499.6 0
0
28
1 0 3 0 0 0 0 2 0 0 10 2
112 403
112 403
1 0 4 0 0 4096 0 3 0 0 11 2
163 412
164 412
1 0 5 0 0 4096 0 4 0 0 12 2
227 421
227 422
1 0 6 0 0 4096 0 5 0 0 13 2
297 431
297 432
1 0 7 0 0 4096 0 6 0 0 27 2
399 397
399 398
0 1 8 0 0 8192 0 0 1 28 0 3
397 343
397 333
416 333
1 1 9 0 0 8320 0 15 7 0 0 3
361 498
361 496
355 496
4 1 2 0 0 12288 0 15 8 0 0 4
415 507
437 507
437 536
394 536
2 1 2 0 0 12416 0 15 8 0 0 4
355 507
345 507
345 536
394 536
7 1 3 0 0 8320 0 17 12 0 0 5
99 322
76 322
76 403
126 403
126 431
0 1 4 0 0 4224 0 0 11 16 0 4
171 323
171 404
164 404
164 431
0 1 5 0 0 4224 0 0 10 20 0 4
245 325
245 422
199 422
199 432
0 1 6 0 0 4224 0 0 9 23 0 3
315 325
315 432
236 432
3 0 10 0 0 8320 0 13 0 0 15 3
171 246
161 246
161 322
2 4 10 0 0 0 0 17 17 0 0 4
147 322
161 322
161 340
147 340
2 7 4 0 0 0 0 13 18 0 0 5
216 255
216 290
171 290
171 323
175 323
0 3 11 0 0 4096 0 0 14 18 0 2
228 249
247 249
0 1 11 0 0 4224 0 0 13 19 0 3
228 323
228 237
216 237
2 4 11 0 0 0 0 18 18 0 0 4
223 323
229 323
229 341
223 341
2 7 5 0 0 0 0 14 19 0 0 5
292 258
292 289
245 289
245 325
252 325
0 1 6 0 0 0 0 0 14 22 0 3
304 325
304 240
292 240
4 0 6 0 0 0 0 19 0 0 23 3
300 343
304 343
304 325
2 7 6 0 0 0 0 19 16 0 0 2
300 325
322 325
3 0 7 0 0 8192 0 19 0 0 26 3
300 334
310 334
310 398
3 0 7 0 0 8192 0 18 0 0 26 3
223 332
235 332
235 398
0 3 7 0 0 4224 0 0 17 27 0 4
373 398
157 398
157 331
147 331
3 3 7 0 0 0 0 15 16 0 0 4
409 498
409 398
370 398
370 334
2 4 8 0 0 4224 0 16 16 0 0 4
370 325
405 325
405 343
370 343
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
