CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 172 63 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5551 0 0
2
44499.9 0
0
13 Logic Switch~
5 276 66 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6986 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 242 66 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8745 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 217 55 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9592 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 139 69 0 1 11
0 23
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8748 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 99 61 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7168 0 0
2
5.90006e-315 0
0
9 Inverter~
13 328 581 0 2 22
0 22 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
631 0 0
2
44499.9 0
0
9 Inverter~
13 341 529 0 2 22
0 23 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9466 0 0
2
44499.9 0
0
9 Inverter~
13 338 475 0 2 22
0 24 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3266 0 0
2
44499.9 0
0
8 3-In OR~
219 681 525 0 4 22
0 21 19 18 10
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 8 0
1 U
7693 0 0
2
5.90006e-315 0
0
8 3-In OR~
219 657 348 0 4 22
0 13 14 12 8
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
3723 0 0
2
5.90006e-315 0
0
5 7415~
219 612 165 0 4 22
0 16 3 28 27
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
3440 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 514 563 0 3 22
0 3 17 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6263 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 431 590 0 3 22
0 5 4 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
4900 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 430 484 0 3 22
0 7 4 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8783 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 434 538 0 3 22
0 6 2 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3221 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 575 377 0 3 22
0 16 9 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3215 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 437 411 0 3 22
0 22 25 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7903 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 435 358 0 3 22
0 23 26 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7121 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 438 300 0 3 22
0 24 11 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4484 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 572 319 0 3 22
0 3 15 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5996 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 514 508 0 3 22
0 16 20 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7804 0 0
2
5.90006e-315 0
0
6 74136~
219 428 235 0 3 22
0 24 4 28
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5523 0 0
2
5.90006e-315 0
0
6 74136~
219 425 162 0 3 22
0 23 2 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3330 0 0
2
5.90006e-315 0
0
6 74136~
219 423 97 0 3 22
0 22 4 16
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U2A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3465 0 0
2
5.90006e-315 0
0
9 Inverter~
13 343 368 0 2 22
0 2 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8396 0 0
2
5.90006e-315 0
0
9 Inverter~
13 368 310 0 2 22
0 4 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3685 0 0
2
5.90006e-315 0
0
9 Inverter~
13 349 421 0 2 22
0 4 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7849 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 675 99 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 735 323 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 746 496 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
5.90006e-315 0
0
47
0 0 2 0 0 8192 0 0 0 29 14 3
348 546
242 546
242 358
1 0 3 0 0 4096 0 21 0 0 3 2
548 310
490 310
1 0 3 0 0 4224 0 13 0 0 41 4
490 554
490 256
571 256
571 165
0 0 4 0 0 4096 0 0 0 28 30 2
275 479
275 592
2 1 5 0 0 4224 0 7 14 0 0 2
349 581
407 581
2 1 6 0 0 4224 0 8 16 0 0 2
362 529
410 529
2 1 7 0 0 4224 0 9 15 0 0 2
359 475
406 475
1 4 8 0 0 8320 0 30 11 0 0 3
735 341
735 348
690 348
2 0 4 0 0 4096 0 25 0 0 30 2
407 106
208 106
2 3 9 0 0 12416 0 17 18 0 0 4
551 386
513 386
513 411
458 411
1 4 10 0 0 8320 0 31 10 0 0 3
746 514
746 525
714 525
0 0 4 0 0 0 0 0 0 28 43 3
275 266
276 266
276 244
1 0 4 0 0 0 0 28 0 0 30 2
334 421
208 421
1 0 2 0 0 8320 0 26 0 0 45 3
328 368
242 368
242 171
1 0 4 0 0 0 0 27 0 0 28 2
353 310
275 310
2 2 11 0 0 8320 0 20 27 0 0 3
414 309
414 310
389 310
3 3 12 0 0 8320 0 11 17 0 0 3
644 357
644 377
596 377
1 3 13 0 0 12416 0 11 21 0 0 4
644 339
623 339
623 319
593 319
3 2 14 0 0 4224 0 19 11 0 0 4
456 358
631 358
631 348
645 348
2 3 15 0 0 4224 0 21 20 0 0 4
548 328
462 328
462 300
459 300
1 0 16 0 0 4096 0 17 0 0 22 2
551 368
468 368
1 0 16 0 0 8320 0 22 0 0 42 3
490 499
468 499
468 97
2 3 17 0 0 4224 0 13 14 0 0 4
490 572
466 572
466 590
452 590
3 3 18 0 0 4224 0 10 13 0 0 6
668 534
591 534
591 577
557 577
557 563
535 563
3 2 19 0 0 12416 0 22 10 0 0 4
535 508
583 508
583 525
669 525
3 2 20 0 0 4224 0 16 22 0 0 4
455 538
476 538
476 517
490 517
3 1 21 0 0 12416 0 15 10 0 0 6
451 484
478 484
478 454
640 454
640 516
668 516
2 0 4 0 0 12416 0 15 0 0 0 4
406 493
406 490
275 490
275 261
2 0 2 0 0 128 0 16 0 0 0 3
410 547
410 546
344 546
2 1 4 0 0 16512 0 14 4 0 0 6
407 599
389 599
389 592
208 592
208 67
217 67
0 1 22 0 0 8192 0 0 7 35 0 3
102 392
102 581
313 581
0 1 23 0 0 4096 0 0 8 36 0 3
141 341
141 529
326 529
0 1 24 0 0 4096 0 0 9 38 0 3
171 244
171 475
323 475
2 2 25 0 0 8320 0 28 18 0 0 3
370 421
370 420
413 420
1 0 22 0 0 8320 0 18 0 0 47 3
413 402
102 402
102 88
1 0 23 0 0 4224 0 19 0 0 46 4
411 349
141 349
141 148
140 148
2 2 26 0 0 8320 0 26 19 0 0 3
364 368
364 367
411 367
1 0 24 0 0 4224 0 20 0 0 44 4
414 291
171 291
171 209
172 209
4 1 27 0 0 8320 0 12 29 0 0 3
633 165
675 165
675 117
3 3 28 0 0 4224 0 12 23 0 0 4
588 174
487 174
487 235
461 235
2 3 3 0 0 0 0 12 24 0 0 4
588 165
481 165
481 162
458 162
3 1 16 0 0 0 0 25 12 0 0 4
456 97
533 97
533 156
588 156
2 1 4 0 0 0 0 23 2 0 0 3
412 244
276 244
276 78
1 1 24 0 0 0 0 1 23 0 0 5
172 75
172 211
353 211
353 226
412 226
2 1 2 0 0 0 0 24 3 0 0 3
409 171
242 171
242 78
1 1 23 0 0 0 0 5 24 0 0 4
139 81
140 81
140 153
409 153
1 1 22 0 0 0 0 6 25 0 0 4
99 73
102 73
102 88
407 88
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
786 513 827 534
794 519 818 534
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
772 343 813 364
780 350 804 365
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
709 135 752 156
718 142 742 157
3 A=B
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
