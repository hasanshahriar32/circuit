CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 502
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.312600 0.500000
176 511 1364 707
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 212 116 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5776 0 0
2
5.90027e-315 0
0
13 Logic Switch~
5 221 290 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7207 0 0
2
5.90027e-315 0
0
9 Inverter~
13 106 170 0 2 22
0 4 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4459 0 0
2
44664.5 0
0
9 Inverter~
13 105 137 0 2 22
0 6 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U9A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3760 0 0
2
44664.5 0
0
5 7422~
219 183 143 0 5 22
0 7 5 9 8 3
0
0 0 624 0
6 74LS22
-21 -28 21 -20
3 U8A
-12 -31 9 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 3 0
1 U
754 0 0
2
44664.5 0
0
5 SCOPE
12 294 135 0 1 11
0 7
0
0 0 57584 270
3 TP5
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9767 0 0
2
44664.5 0
0
5 SCOPE
12 431 134 0 1 11
0 6
0
0 0 57584 270
3 TP4
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7978 0 0
2
44664.5 0
0
5 SCOPE
12 549 135 0 1 11
0 5
0
0 0 57584 270
3 TP3
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3142 0 0
2
44664.5 0
0
5 SCOPE
12 667 135 0 1 11
0 4
0
0 0 57584 270
3 TP2
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3284 0 0
2
44664.5 0
0
5 SCOPE
12 783 145 0 1 11
0 10
0
0 0 57584 270
3 TP1
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
659 0 0
2
44664.5 0
0
7 Pulser~
4 828 221 0 10 12
0 11 2 10 2 0 0 5 5 4
7
0
0 0 4656 180
0
2 V4
-7 -29 7 -21
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 V
3800 0 0
2
44664.4 0
0
2 +V
167 899 157 0 1 3
0 11
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6792 0 0
2
5.90027e-315 0
0
7 Ground~
168 825 265 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 287 77 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 422 78 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 540 77 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7988 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 659 82 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3217 0 0
2
5.90027e-315 0
0
14 Logic Display~
6 775 80 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3965 0 0
2
5.90027e-315 0
0
6 74112~
219 337 255 0 7 32
0 13 12 6 12 3 14 7
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U2B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8239 0 0
2
5.90027e-315 0
0
6 74112~
219 464 255 0 7 32
0 13 12 5 12 3 15 6
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U2A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
828 0 0
2
5.90027e-315 0
0
6 74112~
219 584 255 0 7 32
0 13 12 4 12 3 16 5
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U1B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
6187 0 0
2
5.90027e-315 0
0
6 74112~
219 702 255 0 7 32
0 13 12 10 12 3 17 4
0
0 0 4720 180
5 74112
4 -60 39 -52
3 U1A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
7107 0 0
2
5.90027e-315 0
0
40
5 0 3 0 0 4096 0 5 0 0 37 3
210 143
245 143
245 166
1 1 4 0 0 12416 0 3 17 0 0 6
91 170
27 170
27 23
645 23
645 100
659 100
2 0 5 0 0 12416 0 5 0 0 19 6
159 149
41 149
41 39
517 39
517 99
540 99
1 0 6 0 0 12416 0 4 0 0 20 6
90 137
54 137
54 54
365 54
365 100
422 100
1 1 7 0 0 12416 0 5 14 0 0 4
159 125
133 125
133 95
287 95
2 4 8 0 0 4224 0 3 5 0 0 4
127 170
152 170
152 161
159 161
2 3 9 0 0 4224 0 4 5 0 0 2
126 137
159 137
1 0 7 0 0 0 0 6 0 0 21 2
285 138
287 138
1 0 6 0 0 0 0 7 0 0 20 2
422 137
422 137
1 0 5 0 0 0 0 8 0 0 19 2
540 138
540 138
1 0 4 0 0 0 0 9 0 0 18 2
658 138
659 138
1 0 10 0 0 4096 0 10 0 0 13 2
774 148
775 148
0 1 10 0 0 4224 0 0 18 17 0 2
775 228
775 98
1 0 2 0 0 0 0 13 0 0 15 2
825 259
825 259
4 2 2 0 0 12416 0 11 11 0 0 6
798 219
786 219
786 259
867 259
867 219
858 219
1 1 11 0 0 8320 0 11 12 0 0 3
852 228
899 228
899 166
3 3 10 0 0 0 0 22 11 0 0 2
732 228
804 228
1 0 4 0 0 128 0 17 0 0 38 2
659 100
659 237
1 0 5 0 0 128 0 16 0 0 39 2
540 95
540 237
1 0 6 0 0 128 0 15 0 0 40 2
422 96
422 237
1 7 7 0 0 128 0 14 19 0 0 3
287 95
287 237
313 237
4 0 12 0 0 4096 0 19 0 0 23 2
361 219
388 219
2 0 12 0 0 8192 0 19 0 0 29 3
361 237
388 237
388 116
4 0 12 0 0 0 0 20 0 0 25 2
488 219
512 219
2 0 12 0 0 0 0 20 0 0 29 3
488 237
512 237
512 116
4 0 12 0 0 0 0 21 0 0 27 2
608 219
629 219
2 0 12 0 0 0 0 21 0 0 29 3
608 237
629 237
629 116
4 0 12 0 0 0 0 22 0 0 29 2
726 219
762 219
1 2 12 0 0 4224 0 1 22 0 0 4
224 116
762 116
762 237
726 237
1 0 13 0 0 4096 0 19 0 0 33 2
337 264
337 290
1 0 13 0 0 0 0 20 0 0 33 2
464 264
464 290
1 0 13 0 0 0 0 21 0 0 33 2
584 264
584 290
1 1 13 0 0 4224 0 2 22 0 0 3
233 290
702 290
702 264
5 0 3 0 0 0 0 19 0 0 37 2
337 189
337 166
5 0 3 0 0 0 0 20 0 0 37 2
464 189
464 166
5 0 3 0 0 0 0 21 0 0 37 2
584 189
584 166
0 5 3 0 0 4224 0 0 22 0 0 3
230 166
702 166
702 189
3 7 4 0 0 0 0 21 22 0 0 4
614 228
646 228
646 237
678 237
3 7 5 0 0 0 0 20 21 0 0 4
494 228
529 228
529 237
560 237
3 7 6 0 0 0 0 19 20 0 0 4
367 228
402 228
402 237
440 237
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
