CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 168 217 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44664.5 0
0
13 Logic Switch~
5 561 133 0 1 11
0 18
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44664.5 1
0
13 Logic Switch~
5 560 328 0 1 11
0 19
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
44664.5 2
0
13 Logic Switch~
5 702 323 0 1 11
0 16
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44664.5 3
0
13 Logic Switch~
5 703 128 0 1 11
0 15
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44664.5 4
0
13 Logic Switch~
5 422 140 0 1 11
0 21
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
44664.5 5
0
13 Logic Switch~
5 421 335 0 1 11
0 22
0
0 0 21360 90
2 0V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44664.5 6
0
13 Logic Switch~
5 279 340 0 1 11
0 25
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
44664.5 7
0
13 Logic Switch~
5 280 145 0 1 11
0 24
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
44664.5 8
0
9 Inverter~
13 505 230 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
972 0 0
2
44664.5 9
0
9 Inverter~
13 652 225 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3472 0 0
2
44664.5 10
0
9 Inverter~
13 368 236 0 2 22
0 9 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9998 0 0
2
44664.5 11
0
9 Inverter~
13 200 241 0 2 22
0 11 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3536 0 0
2
44664.5 12
0
14 Logic Display~
6 203 274 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90027e-315 0
0
2 +V
167 81 286 0 1 3
0 12
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
5.90027e-315 5.26354e-315
0
7 Ground~
168 90 370 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3670 0 0
2
5.90027e-315 5.30499e-315
0
7 Pulser~
4 151 321 0 10 12
0 12 2 3 2 0 0 10 10 3
8
0
0 0 4656 0
0
3 V10
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 V
5616 0 0
2
44664.5 13
0
5 4027~
219 561 246 0 7 32
0 18 7 3 6 19 17 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 2 0
1 U
9323 0 0
2
44664.5 14
0
14 Logic Display~
6 609 165 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
44664.5 15
0
14 Logic Display~
6 610 282 0 1 2
10 17
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
44664.5 16
0
14 Logic Display~
6 752 277 0 1 2
10 13
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
44664.5 17
0
14 Logic Display~
6 751 160 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
44664.5 18
0
5 4027~
219 703 241 0 7 32
0 15 5 3 4 16 13 14
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
7876 0 0
2
44664.5 19
0
5 4027~
219 422 253 0 7 32
0 21 9 3 8 22 20 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 1 0
1 U
6369 0 0
2
44664.5 20
0
14 Logic Display~
6 470 172 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
44664.5 21
0
14 Logic Display~
6 471 289 0 1 2
10 20
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
44664.5 22
0
14 Logic Display~
6 329 294 0 1 2
10 23
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
44664.5 23
0
14 Logic Display~
6 328 177 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
44664.5 24
0
5 4027~
219 280 258 0 7 32
0 24 11 3 10 25 23 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 1 0
1 U
961 0 0
2
44664.5 25
0
36
0 3 3 0 0 8320 0 0 23 12 0 4
519 382
673 382
673 214
679 214
2 4 4 0 0 8320 0 11 23 0 0 3
673 225
673 223
679 223
1 0 5 0 0 8192 0 11 0 0 18 3
637 225
633 225
633 205
2 4 6 0 0 12416 0 10 18 0 0 4
526 230
531 230
531 228
537 228
1 0 7 0 0 8192 0 10 0 0 19 3
490 230
486 230
486 210
2 4 8 0 0 8320 0 12 24 0 0 3
389 236
389 235
398 235
1 0 9 0 0 8192 0 12 0 0 20 3
353 236
349 236
349 217
2 4 10 0 0 4224 0 13 29 0 0 4
221 241
248 241
248 240
256 240
0 1 11 0 0 12288 0 0 13 17 0 5
186 217
186 227
177 227
177 241
185 241
3 0 3 0 0 0 0 29 0 0 13 5
256 231
237 231
237 382
203 382
203 312
3 0 3 0 0 0 0 24 0 0 10 4
398 226
374 226
374 382
237 382
3 0 3 0 0 0 0 18 0 0 11 4
537 219
519 219
519 382
374 382
3 1 3 0 0 0 0 17 14 0 0 3
175 312
203 312
203 292
1 1 12 0 0 8320 0 15 17 0 0 3
81 295
81 312
127 312
2 0 2 0 0 8192 0 17 0 0 16 3
121 321
91 321
91 356
4 1 2 0 0 12416 0 17 16 0 0 5
181 321
185 321
185 356
90 356
90 364
1 2 11 0 0 4224 0 1 29 0 0 4
180 217
248 217
248 222
256 222
0 2 5 0 0 8320 0 0 23 26 0 3
609 210
609 205
679 205
0 2 7 0 0 8320 0 0 18 30 0 3
469 217
469 210
537 210
0 2 9 0 0 8320 0 0 24 34 0 3
328 222
328 217
398 217
6 1 13 0 0 8320 0 23 21 0 0 3
733 223
752 223
752 263
7 1 14 0 0 8320 0 23 22 0 0 3
727 205
751 205
751 178
1 1 15 0 0 4224 0 23 5 0 0 2
703 184
703 140
1 5 16 0 0 4224 0 4 23 0 0 2
703 310
703 247
6 1 17 0 0 8320 0 18 20 0 0 3
591 228
610 228
610 268
7 1 5 0 0 0 0 18 19 0 0 3
585 210
609 210
609 183
1 1 18 0 0 4224 0 18 2 0 0 2
561 189
561 145
1 5 19 0 0 4224 0 3 18 0 0 2
561 315
561 252
6 1 20 0 0 8320 0 24 26 0 0 3
452 235
471 235
471 275
7 1 7 0 0 0 0 24 25 0 0 3
446 217
470 217
470 190
1 1 21 0 0 4224 0 24 6 0 0 2
422 196
422 152
1 5 22 0 0 4224 0 7 24 0 0 2
422 322
422 259
6 1 23 0 0 8320 0 29 27 0 0 3
310 240
329 240
329 280
7 1 9 0 0 0 0 29 28 0 0 3
304 222
328 222
328 195
1 1 24 0 0 4224 0 29 9 0 0 2
280 201
280 157
1 5 25 0 0 4224 0 8 29 0 0 2
280 327
280 264
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
774 66 827 90
784 74 816 90
4 SISO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
493 78 546 102
503 86 535 102
4 SISO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
