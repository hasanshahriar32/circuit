CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 554 363 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44500.1 0
0
13 Logic Switch~
5 510 353 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44500.1 0
0
13 Logic Switch~
5 552 300 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
44500.1 0
0
13 Logic Switch~
5 510 277 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
44500.1 0
0
13 Logic Switch~
5 549 225 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
44500.1 0
0
13 Logic Switch~
5 503 213 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44500.1 0
0
13 Logic Switch~
5 543 146 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
44500.1 0
0
13 Logic Switch~
5 496 127 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
44500.1 0
0
13 Logic Switch~
5 171 302 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 197 248 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 161 221 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 204 169 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90006e-315 0
0
13 Logic Switch~
5 164 142 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 730 330 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44500.1 0
0
14 Logic Display~
6 730 264 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
44500.1 0
0
14 Logic Display~
6 732 188 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
44500.1 0
0
14 Logic Display~
6 730 101 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44500.1 0
0
6 74266~
219 617 358 0 3 22
0 7 6 5
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
9323 0 0
2
44500.1 0
0
6 74136~
219 615 289 0 3 22
0 9 8 4
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
317 0 0
2
44500.1 0
0
9 2-In NOR~
219 614 219 0 3 22
0 11 10 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3108 0 0
2
44500.1 0
0
10 2-In NAND~
219 624 135 0 3 22
0 13 12 2
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4299 0 0
2
44500.1 0
0
14 Logic Display~
6 414 281 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 414 216 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.90006e-315 0
0
14 Logic Display~
6 415 143 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.90006e-315 0
0
9 Inverter~
13 325 302 0 2 22
0 17 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9172 0 0
2
5.90006e-315 0
0
8 2-In OR~
219 321 240 0 3 22
0 19 18 15
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7100 0 0
2
5.90006e-315 0
0
9 2-In AND~
219 331 165 0 3 22
0 21 20 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3820 0 0
2
5.90006e-315 0
0
20
3 1 2 0 0 4224 0 21 17 0 0 3
651 135
730 135
730 119
3 1 3 0 0 4224 0 20 16 0 0 3
653 219
732 219
732 206
3 1 4 0 0 4224 0 19 15 0 0 3
648 289
730 289
730 282
3 1 5 0 0 4224 0 18 14 0 0 3
656 358
730 358
730 348
2 1 6 0 0 4224 0 18 1 0 0 4
601 367
575 367
575 363
566 363
1 1 7 0 0 4224 0 18 2 0 0 4
601 349
531 349
531 353
522 353
1 2 8 0 0 4224 0 3 19 0 0 4
564 300
591 300
591 298
599 298
1 1 9 0 0 4224 0 19 4 0 0 4
599 280
531 280
531 277
522 277
2 1 10 0 0 4224 0 20 5 0 0 4
601 228
570 228
570 225
561 225
1 1 11 0 0 4224 0 20 6 0 0 4
601 210
524 210
524 213
515 213
2 1 12 0 0 4224 0 21 7 0 0 4
600 144
564 144
564 146
555 146
1 1 13 0 0 4224 0 21 8 0 0 4
600 126
517 126
517 127
508 127
3 1 14 0 0 4224 0 27 24 0 0 3
352 165
415 165
415 161
3 1 15 0 0 4224 0 26 23 0 0 3
354 240
414 240
414 234
2 1 16 0 0 4224 0 25 22 0 0 3
346 302
414 302
414 299
1 1 17 0 0 4224 0 9 25 0 0 2
183 302
310 302
1 2 18 0 0 4224 0 10 26 0 0 4
209 248
300 248
300 249
308 249
1 1 19 0 0 4224 0 11 26 0 0 4
173 221
300 221
300 231
308 231
1 2 20 0 0 4224 0 12 27 0 0 4
216 169
299 169
299 174
307 174
1 1 21 0 0 4224 0 13 27 0 0 4
176 142
299 142
299 156
307 156
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
