CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 440 1364 717
9437202 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 123 109 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -32 8 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
44500.2 0
0
13 Logic Switch~
5 284 118 0 1 11
0 3
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6369 0 0
2
44500.2 0
0
13 Logic Switch~
5 232 112 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
44500.2 2
0
13 Logic Switch~
5 175 126 0 1 11
0 4
0
0 0 21360 270
2 0V
-7 -21 7 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7100 0 0
2
44500.2 3
0
9 2-In AND~
219 325 488 0 3 22
0 4 3 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3820 0 0
2
44500.2 0
0
9 2-In AND~
219 325 446 0 3 22
0 4 2 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7678 0 0
2
44500.2 0
0
8 3-In OR~
219 435 439 0 4 22
0 5 6 7 16
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 6 0
1 U
961 0 0
2
44500.2 0
0
8 3-In OR~
219 399 305 0 4 22
0 10 9 8 15
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
3178 0 0
2
44500.2 0
0
5 7415~
219 340 365 0 4 22
0 4 12 11 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
3409 0 0
2
44500.2 0
0
9 2-In AND~
219 343 318 0 3 22
0 13 3 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3951 0 0
2
44500.2 0
0
9 2-In AND~
219 343 263 0 3 22
0 13 2 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8885 0 0
2
44500.2 0
0
9 Inverter~
13 247 169 0 2 22
0 2 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3780 0 0
2
44500.2 0
0
9 Inverter~
13 190 161 0 2 22
0 4 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9265 0 0
2
44500.2 0
0
6 74266~
219 385 196 0 3 22
0 2 3 14
0
0 0 624 0
7 74LS266
-24 -24 25 -16
3 U2B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9442 0 0
2
44500.2 4
0
14 Logic Display~
6 553 420 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
44500.2 5
0
14 Logic Display~
6 545 255 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
44500.2 6
0
14 Logic Display~
6 546 186 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
44500.2 7
0
14 Logic Display~
6 546 101 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
44500.2 8
0
9 Inverter~
13 299 148 0 2 22
0 3 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7168 0 0
2
44500.2 13
0
32
1 0 2 0 0 4096 0 14 0 0 25 2
369 187
232 187
2 0 3 0 0 4096 0 5 0 0 22 2
301 497
284 497
1 0 4 0 0 4096 0 5 0 0 28 2
301 479
175 479
2 0 2 0 0 0 0 6 0 0 25 2
301 455
232 455
1 0 4 0 0 0 0 6 0 0 28 2
301 437
175 437
1 0 5 0 0 4096 0 7 0 0 21 2
422 430
123 430
2 3 6 0 0 4224 0 7 6 0 0 4
423 439
362 439
362 446
346 446
3 3 7 0 0 12416 0 5 7 0 0 4
346 488
368 488
368 448
422 448
3 4 8 0 0 8320 0 8 9 0 0 4
386 314
374 314
374 365
361 365
2 3 9 0 0 4224 0 8 10 0 0 4
387 305
370 305
370 318
364 318
1 3 10 0 0 8320 0 8 11 0 0 4
386 296
370 296
370 263
364 263
3 0 11 0 0 8192 0 9 0 0 32 5
316 374
301 374
301 172
328 172
328 148
2 0 12 0 0 4096 0 9 0 0 24 2
316 365
268 365
1 0 4 0 0 4096 0 9 0 0 28 2
316 356
175 356
2 0 3 0 0 4096 0 10 0 0 22 2
319 327
284 327
1 0 13 0 0 4096 0 10 0 0 26 2
319 309
211 309
2 0 2 0 0 0 0 11 0 0 25 2
319 272
232 272
1 0 13 0 0 0 0 11 0 0 26 2
319 254
211 254
2 0 3 0 0 4096 0 14 0 0 22 2
369 205
284 205
1 0 3 0 0 0 0 19 0 0 22 2
284 148
284 148
1 0 5 0 0 4224 0 1 0 0 0 2
123 121
123 654
1 0 3 0 0 4224 0 2 0 0 0 2
284 130
284 712
1 0 2 0 0 0 0 12 0 0 25 2
232 169
232 169
2 0 12 0 0 4224 0 12 0 0 0 4
268 169
268 673
276 673
276 688
1 0 2 0 0 4224 0 3 0 0 0 2
232 124
232 663
2 0 13 0 0 4224 0 13 0 0 0 2
211 161
211 603
1 0 4 0 0 0 0 13 0 0 28 2
175 161
175 161
1 0 4 0 0 4224 0 4 0 0 0 2
175 138
175 606
1 3 14 0 0 8320 0 17 14 0 0 4
546 204
546 212
424 212
424 196
4 1 15 0 0 4224 0 8 16 0 0 3
432 305
545 305
545 273
1 4 16 0 0 8320 0 15 7 0 0 5
553 438
553 443
477 443
477 439
468 439
1 2 11 0 0 12416 0 18 19 0 0 4
546 119
531 119
531 148
320 148
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
599 428 626 449
608 435 616 450
1 W
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
589 288 616 309
598 295 606 310
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
592 193 617 214
600 199 608 214
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
573 113 600 134
582 119 590 134
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
270 55 297 76
279 62 287 77
1 D
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
225 41 250 62
233 48 241 63
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
167 56 192 77
175 63 183 78
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
108 51 135 72
117 58 125 73
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
