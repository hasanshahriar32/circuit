CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 660 30 90 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 365 121 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8323 0 0
2
5.90003e-315 0
0
13 Logic Switch~
5 208 125 0 1 11
0 13
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3984 0 0
2
5.90003e-315 5.26354e-315
0
13 Logic Switch~
5 50 129 0 1 11
0 14
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7622 0 0
2
5.90003e-315 0
0
14 Logic Display~
6 744 1082 0 1 2
10 3
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L10
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
816 0 0
2
44500 0
0
8 4-In OR~
219 763 1030 0 5 22
0 2 4 5 6 3
0
0 0 624 270
4 4072
-14 -24 14 -16
3 U5B
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
4656 0 0
2
44500 0
0
8 4-In OR~
219 710 1034 0 5 22
0 2 8 9 10 7
0
0 0 624 270
4 4072
-14 -24 14 -16
3 U5A
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
6356 0 0
2
44500 0
0
14 Logic Display~
6 688 1086 0 1 2
10 7
0
0 0 53856 90
6 100MEG
3 -16 45 -8
2 L9
-9 -15 5 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7479 0 0
2
44500 0
0
5 7415~
219 651 530 0 4 22
0 14 15 12 8
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
5690 0 0
2
5.90003e-315 5.37752e-315
0
14 Logic Display~
6 786 522 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5617 0 0
2
5.90003e-315 5.36716e-315
0
14 Logic Display~
6 787 601 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3903 0 0
2
5.90003e-315 5.3568e-315
0
5 7415~
219 652 609 0 4 22
0 14 15 11 5
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
4452 0 0
2
5.90003e-315 5.34643e-315
0
5 7415~
219 651 773 0 4 22
0 14 13 11 2
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
6282 0 0
2
5.90003e-315 5.32571e-315
0
14 Logic Display~
6 786 765 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7187 0 0
2
5.90003e-315 5.30499e-315
0
14 Logic Display~
6 785 686 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6866 0 0
2
5.90003e-315 5.26354e-315
0
5 7415~
219 650 694 0 4 22
0 14 13 12 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 2 0
1 U
7670 0 0
2
5.90003e-315 0
0
5 7415~
219 650 380 0 4 22
0 16 13 12 9
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 2 0
1 U
951 0 0
2
5.90003e-315 5.32571e-315
0
14 Logic Display~
6 785 372 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9536 0 0
2
5.90003e-315 5.30499e-315
0
14 Logic Display~
6 786 451 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5495 0 0
2
5.90003e-315 5.26354e-315
0
5 7415~
219 651 459 0 4 22
0 16 13 11 6
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 2 0
1 U
8152 0 0
2
5.90003e-315 0
0
5 7415~
219 652 295 0 4 22
0 16 15 11 10
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 1 0
1 U
6223 0 0
2
5.90003e-315 5.26354e-315
0
14 Logic Display~
6 787 287 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5441 0 0
2
5.90003e-315 0
0
14 Logic Display~
6 786 208 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3189 0 0
2
5.90003e-315 0
0
9 Inverter~
13 423 165 0 2 22
0 11 12
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8460 0 0
2
5.90003e-315 5.26354e-315
0
9 Inverter~
13 266 169 0 2 22
0 13 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5179 0 0
2
5.90003e-315 0
0
9 Inverter~
13 108 175 0 2 22
0 14 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U4A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3593 0 0
2
5.90003e-315 0
0
5 7415~
219 651 216 0 4 22
0 16 15 12 17
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 1 0
1 U
3928 0 0
2
5.90003e-315 0
0
54
1 0 2 0 0 4224 0 6 0 0 39 2
726 1014
726 773
5 1 3 0 0 12416 0 5 4 0 0 4
766 1060
766 1067
759 1067
759 1085
1 0 2 0 0 0 0 5 0 0 39 2
779 1010
779 791
2 0 4 0 0 4224 0 5 0 0 40 2
770 1010
770 694
3 0 5 0 0 4224 0 5 0 0 41 2
761 1010
761 609
4 0 6 0 0 4224 0 5 0 0 43 2
752 1010
752 459
5 1 7 0 0 4224 0 6 7 0 0 3
713 1064
713 1089
703 1089
2 0 8 0 0 4096 0 6 0 0 11 2
717 1014
717 1010
3 0 9 0 0 4096 0 6 0 0 12 2
708 1014
708 1010
4 0 10 0 0 4096 0 6 0 0 13 2
699 1014
699 1010
0 0 8 0 0 4224 0 0 0 0 42 2
717 1016
717 530
0 0 9 0 0 4224 0 0 0 0 44 2
708 1016
708 380
0 0 10 0 0 4224 0 0 0 45 0 4
680 295
680 980
699 980
699 1014
0 3 11 0 0 4096 0 0 12 48 0 2
365 782
627 782
0 3 12 0 0 4096 0 0 15 47 0 2
426 703
626 703
0 2 13 0 0 4096 0 0 12 51 0 2
208 773
627 773
0 2 13 0 0 0 0 0 15 51 0 2
208 694
626 694
0 1 14 0 0 4096 0 0 8 22 0 2
50 521
627 521
0 1 14 0 0 4096 0 0 11 22 0 2
50 600
628 600
0 1 14 0 0 0 0 0 15 22 0 2
50 685
626 685
0 1 14 0 0 0 0 0 12 22 0 2
50 764
627 764
0 0 14 0 0 4224 0 0 0 54 0 2
50 149
50 899
0 3 11 0 0 4096 0 0 11 48 0 2
365 618
628 618
0 2 15 0 0 4096 0 0 11 50 0 2
269 609
628 609
0 3 12 0 0 4096 0 0 8 47 0 2
426 539
627 539
0 2 15 0 0 0 0 0 8 50 0 2
269 530
627 530
0 3 11 0 0 0 0 0 19 48 0 2
365 468
627 468
0 2 13 0 0 0 0 0 19 51 0 2
208 459
627 459
0 1 16 0 0 4096 0 0 19 53 0 2
111 450
627 450
0 3 12 0 0 0 0 0 16 47 0 2
426 389
626 389
0 2 13 0 0 0 0 0 16 51 0 2
208 380
626 380
0 1 16 0 0 0 0 0 16 53 0 2
111 371
626 371
0 3 11 0 0 0 0 0 20 48 0 2
365 304
628 304
0 2 15 0 0 0 0 0 20 50 0 2
269 295
628 295
0 1 16 0 0 4096 0 0 20 53 0 2
111 286
628 286
0 3 12 0 0 0 0 0 26 47 0 2
426 225
627 225
0 2 15 0 0 0 0 0 26 50 0 2
269 216
627 216
0 1 16 0 0 0 0 0 26 53 0 2
111 207
627 207
4 1 2 0 0 128 0 12 13 0 0 5
672 773
774 773
774 791
786 791
786 783
4 1 4 0 0 128 0 15 14 0 0 5
671 694
773 694
773 712
785 712
785 704
4 1 5 0 0 128 0 11 10 0 0 5
673 609
775 609
775 627
787 627
787 619
4 1 8 0 0 128 0 8 9 0 0 5
672 530
774 530
774 548
786 548
786 540
4 1 6 0 0 128 0 19 18 0 0 5
672 459
774 459
774 477
786 477
786 469
4 1 9 0 0 128 0 16 17 0 0 5
671 380
773 380
773 398
785 398
785 390
4 1 10 0 0 128 0 20 21 0 0 5
673 295
775 295
775 313
787 313
787 305
4 1 17 0 0 4224 0 26 22 0 0 5
672 216
774 216
774 234
786 234
786 226
2 0 12 0 0 4224 0 23 0 0 0 2
426 183
426 830
0 0 11 0 0 4224 0 0 0 49 0 2
365 141
365 896
1 1 11 0 0 0 0 1 23 0 0 4
365 133
365 141
426 141
426 147
2 0 15 0 0 4224 0 24 0 0 0 2
269 187
269 885
0 0 13 0 0 4224 0 0 0 52 0 2
208 145
208 894
1 1 13 0 0 0 0 2 24 0 0 4
208 137
208 145
269 145
269 151
2 0 16 0 0 4224 0 25 0 0 0 2
111 193
111 907
1 1 14 0 0 0 0 3 25 0 0 4
50 141
50 149
111 149
111 157
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
742 1099 771 1123
753 1108 759 1124
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
676 1100 707 1124
688 1109 694 1125
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
34 72 63 96
44 80 52 96
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
192 68 221 92
202 76 210 92
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
349 64 378 88
359 72 367 88
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 194 823 218
796 202 812 218
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
787 273 824 297
797 281 813 297
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 358 822 382
795 366 811 382
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 437 823 461
796 445 812 461
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 508 823 532
796 516 812 532
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
787 587 824 611
797 595 813 611
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 672 822 696
795 680 811 696
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 751 823 775
796 759 812 775
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
562 65 639 89
572 73 628 89
7 Decoder
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
