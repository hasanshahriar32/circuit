CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 10
176 80 1364 513
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.295133 0.500000
176 522 1364 707
76546066 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 82 173 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44663.4 0
0
5 SCOPE
12 219 279 0 1 11
0 3
0
0 0 57568 0
3 CLK
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
391 0 0
2
44663.4 1
0
5 SCOPE
12 240 172 0 1 11
0 4
0
0 0 57568 0
2 Qa
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3124 0 0
2
44663.4 2
0
5 SCOPE
12 364 157 0 1 11
0 5
0
0 0 57568 0
2 Qb
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3421 0 0
2
44663.4 3
0
5 SCOPE
12 469 161 0 1 11
0 6
0
0 0 57568 0
2 Qc
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8157 0 0
2
44663.4 4
0
14 Logic Display~
6 674 165 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
44663.4 5
0
14 Logic Display~
6 540 137 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
44663.4 6
0
14 Logic Display~
6 431 149 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
44663.4 7
0
14 Logic Display~
6 176 273 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
44663.4 8
0
14 Logic Display~
6 328 160 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
44663.4 9
0
14 Logic Display~
6 214 163 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
44663.4 10
0
5 SCOPE
12 569 168 0 1 11
0 7
0
0 0 57568 0
2 Qd
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9998 0 0
2
44663.4 11
0
5 SCOPE
12 702 168 0 1 11
0 8
0
0 0 57568 0
2 Qe
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3536 0 0
2
44663.4 12
0
7 Ground~
168 117 356 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
44663.4 13
0
2 +V
167 40 273 0 1 3
0 13
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3835 0 0
2
44663.4 14
0
7 Pulser~
4 113 310 0 10 12
0 13 2 3 2 0 0 5 5 2
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 V
3670 0 0
2
44663.4 15
0
9 2-In AND~
219 590 92 0 3 22
0 11 7 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5616 0 0
2
44663.4 16
0
9 2-In AND~
219 495 78 0 3 22
0 12 6 11
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9323 0 0
2
44663.4 17
0
9 2-In AND~
219 357 101 0 3 22
0 4 5 12
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
317 0 0
2
44663.4 18
0
5 4027~
219 625 244 0 7 32
0 14 10 3 15 16 17 8
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U3A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
3108 0 0
2
44663.4 19
0
5 4027~
219 516 247 0 7 32
0 18 11 3 19 20 21 7
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
4299 0 0
2
44663.4 20
0
5 4027~
219 417 247 0 7 32
0 22 12 3 23 24 25 6
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9672 0 0
2
44663.4 21
0
5 4027~
219 309 246 0 7 32
0 26 4 3 27 28 29 5
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7876 0 0
2
44663.4 22
0
5 4027~
219 182 247 0 7 32
0 30 9 3 31 32 33 4
0
0 0 4704 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6369 0 0
2
44663.4 23
0
32
1 0 3 0 0 4096 0 2 0 0 29 3
219 291
219 297
221 297
1 0 4 0 0 4096 0 3 0 0 32 2
240 184
240 211
1 0 5 0 0 4096 0 4 0 0 22 2
364 169
343 169
1 0 6 0 0 4096 0 5 0 0 19 2
469 173
441 173
1 0 7 0 0 4096 0 12 0 0 16 2
569 180
548 180
1 0 8 0 0 4096 0 6 0 0 14 2
674 183
702 183
1 0 7 0 0 0 0 7 0 0 16 3
540 155
540 165
548 165
1 0 6 0 0 0 0 8 0 0 19 2
431 167
441 167
1 0 5 0 0 0 0 10 0 0 22 2
328 178
343 178
1 0 4 0 0 4096 0 11 0 0 32 2
214 181
214 211
0 0 3 0 0 4096 0 0 0 29 29 2
165 297
187 297
1 0 3 0 0 0 0 9 0 0 29 2
176 291
176 297
1 2 9 0 0 4224 0 1 24 0 0 4
94 173
150 173
150 211
158 211
7 1 8 0 0 4224 0 20 13 0 0 3
649 208
702 208
702 180
3 2 10 0 0 8320 0 17 20 0 0 6
611 92
615 92
615 183
596 183
596 208
601 208
2 7 7 0 0 8320 0 17 21 0 0 6
566 101
548 101
548 186
554 186
554 211
540 211
0 1 11 0 0 8192 0 0 17 18 0 3
520 78
520 83
566 83
3 2 11 0 0 8320 0 18 21 0 0 6
516 78
520 78
520 185
484 185
484 211
492 211
7 2 6 0 0 4224 0 22 18 0 0 5
441 211
441 125
464 125
464 87
471 87
0 1 12 0 0 4096 0 0 18 21 0 4
385 101
441 101
441 69
471 69
3 2 12 0 0 8320 0 19 22 0 0 4
378 101
385 101
385 211
393 211
7 2 5 0 0 8320 0 23 19 0 0 6
333 210
343 210
343 120
328 120
328 110
333 110
0 1 4 0 0 4224 0 0 19 32 0 3
260 211
260 92
333 92
1 0 2 0 0 4096 0 14 0 0 25 2
117 350
117 337
2 4 2 0 0 12416 0 16 16 0 0 7
83 310
59 310
59 337
156 337
156 313
143 313
143 310
0 3 3 0 0 4224 0 0 20 27 0 4
472 293
595 293
595 217
601 217
0 3 3 0 0 0 0 0 21 28 0 5
376 293
473 293
473 223
492 223
492 220
0 3 3 0 0 0 0 0 22 29 0 4
263 297
376 297
376 220
393 220
0 3 3 0 0 0 0 0 23 30 0 5
150 297
264 297
264 222
285 222
285 219
3 3 3 0 0 0 0 16 24 0 0 4
137 301
150 301
150 220
158 220
1 1 13 0 0 8320 0 15 16 0 0 3
40 282
40 301
89 301
7 2 4 0 0 0 0 24 23 0 0 4
206 211
277 211
277 210
285 210
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
